VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO tdc_64
  CLASS BLOCK ;
  ORIGIN 1.525 35.545 ;
  FOREIGN tdc_64 -1.525 -35.545 ;
  SIZE 956.41 BY 37.77 ;
  SYMMETRY X Y R90 ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT -0.7 -0.35 -0.37 -0.02 ;
    END
  END a
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -1.52 -32.12 954.88 -31.8 ;
        RECT 953.875 -32.125 954.205 -31.795 ;
        RECT 952.515 -32.125 952.845 -31.795 ;
        RECT 951.155 -32.125 951.485 -31.795 ;
        RECT 949.795 -32.125 950.125 -31.795 ;
        RECT 947.075 -32.125 947.405 -31.795 ;
        RECT 945.715 -32.125 946.045 -31.795 ;
        RECT 944.355 -32.125 944.685 -31.795 ;
        RECT 942.995 -32.125 943.325 -31.795 ;
        RECT 941.635 -32.125 941.965 -31.795 ;
        RECT 940.275 -32.125 940.605 -31.795 ;
        RECT 938.915 -32.125 939.245 -31.795 ;
        RECT 937.555 -32.125 937.885 -31.795 ;
        RECT 936.195 -32.125 936.525 -31.795 ;
        RECT 932.115 -32.125 932.445 -31.795 ;
        RECT 928.035 -32.125 928.365 -31.795 ;
        RECT 926.675 -32.125 927.005 -31.795 ;
        RECT 925.315 -32.125 925.645 -31.795 ;
        RECT 923.955 -32.125 924.285 -31.795 ;
        RECT 922.595 -32.125 922.925 -31.795 ;
        RECT 921.235 -32.125 921.565 -31.795 ;
        RECT 917.155 -32.125 917.485 -31.795 ;
        RECT 913.075 -32.125 913.405 -31.795 ;
        RECT 911.715 -32.125 912.045 -31.795 ;
        RECT 910.355 -32.125 910.685 -31.795 ;
        RECT 908.995 -32.125 909.325 -31.795 ;
        RECT 907.635 -32.125 907.965 -31.795 ;
        RECT 906.275 -32.125 906.605 -31.795 ;
        RECT 902.195 -32.125 902.525 -31.795 ;
        RECT 900.835 -32.125 901.165 -31.795 ;
        RECT 898.115 -32.125 898.445 -31.795 ;
        RECT 896.755 -32.125 897.085 -31.795 ;
        RECT 895.395 -32.125 895.725 -31.795 ;
        RECT 894.035 -32.125 894.365 -31.795 ;
        RECT 892.675 -32.125 893.005 -31.795 ;
        RECT 891.315 -32.125 891.645 -31.795 ;
        RECT 885.875 -32.125 886.205 -31.795 ;
        RECT 883.155 -32.125 883.485 -31.795 ;
        RECT 881.795 -32.125 882.125 -31.795 ;
        RECT 880.435 -32.125 880.765 -31.795 ;
        RECT 879.075 -32.125 879.405 -31.795 ;
        RECT 877.715 -32.125 878.045 -31.795 ;
        RECT 876.355 -32.125 876.685 -31.795 ;
        RECT 870.915 -32.125 871.245 -31.795 ;
        RECT 868.195 -32.125 868.525 -31.795 ;
        RECT 866.835 -32.125 867.165 -31.795 ;
        RECT 865.475 -32.125 865.805 -31.795 ;
        RECT 864.115 -32.125 864.445 -31.795 ;
        RECT 862.755 -32.125 863.085 -31.795 ;
        RECT 861.395 -32.125 861.725 -31.795 ;
        RECT 855.955 -32.125 856.285 -31.795 ;
        RECT 853.235 -32.125 853.565 -31.795 ;
        RECT 851.875 -32.125 852.205 -31.795 ;
        RECT 850.515 -32.125 850.845 -31.795 ;
        RECT 849.155 -32.125 849.485 -31.795 ;
        RECT 847.795 -32.125 848.125 -31.795 ;
        RECT 846.435 -32.125 846.765 -31.795 ;
        RECT 843.715 -32.125 844.045 -31.795 ;
        RECT 840.995 -32.125 841.325 -31.795 ;
        RECT 838.275 -32.125 838.605 -31.795 ;
        RECT 836.915 -32.125 837.245 -31.795 ;
        RECT 835.555 -32.125 835.885 -31.795 ;
        RECT 834.195 -32.125 834.525 -31.795 ;
        RECT 832.835 -32.125 833.165 -31.795 ;
        RECT 831.475 -32.125 831.805 -31.795 ;
        RECT 828.755 -32.125 829.085 -31.795 ;
        RECT 826.035 -32.125 826.365 -31.795 ;
        RECT 823.315 -32.125 823.645 -31.795 ;
        RECT 821.955 -32.125 822.285 -31.795 ;
        RECT 820.595 -32.125 820.925 -31.795 ;
        RECT 819.235 -32.125 819.565 -31.795 ;
        RECT 817.875 -32.125 818.205 -31.795 ;
        RECT 816.515 -32.125 816.845 -31.795 ;
        RECT 813.795 -32.125 814.125 -31.795 ;
        RECT 811.075 -32.125 811.405 -31.795 ;
        RECT 808.355 -32.125 808.685 -31.795 ;
        RECT 806.995 -32.125 807.325 -31.795 ;
        RECT 805.635 -32.125 805.965 -31.795 ;
        RECT 804.275 -32.125 804.605 -31.795 ;
        RECT 802.915 -32.125 803.245 -31.795 ;
        RECT 801.555 -32.125 801.885 -31.795 ;
        RECT 798.835 -32.125 799.165 -31.795 ;
        RECT 796.115 -32.125 796.445 -31.795 ;
        RECT 793.395 -32.125 793.725 -31.795 ;
        RECT 792.035 -32.125 792.365 -31.795 ;
        RECT 790.675 -32.125 791.005 -31.795 ;
        RECT 789.315 -32.125 789.645 -31.795 ;
        RECT 787.955 -32.125 788.285 -31.795 ;
        RECT 786.595 -32.125 786.925 -31.795 ;
        RECT 783.875 -32.125 784.205 -31.795 ;
        RECT 781.155 -32.125 781.485 -31.795 ;
        RECT 778.435 -32.125 778.765 -31.795 ;
        RECT 777.075 -32.125 777.405 -31.795 ;
        RECT 775.715 -32.125 776.045 -31.795 ;
        RECT 774.355 -32.125 774.685 -31.795 ;
        RECT 772.995 -32.125 773.325 -31.795 ;
        RECT 771.635 -32.125 771.965 -31.795 ;
        RECT 768.915 -32.125 769.245 -31.795 ;
        RECT 766.195 -32.125 766.525 -31.795 ;
        RECT 763.475 -32.125 763.805 -31.795 ;
        RECT 762.115 -32.125 762.445 -31.795 ;
        RECT 760.755 -32.125 761.085 -31.795 ;
        RECT 759.395 -32.125 759.725 -31.795 ;
        RECT 758.035 -32.125 758.365 -31.795 ;
        RECT 756.675 -32.125 757.005 -31.795 ;
        RECT 753.955 -32.125 754.285 -31.795 ;
        RECT 751.235 -32.125 751.565 -31.795 ;
        RECT 748.515 -32.125 748.845 -31.795 ;
        RECT 747.155 -32.125 747.485 -31.795 ;
        RECT 745.795 -32.125 746.125 -31.795 ;
        RECT 744.435 -32.125 744.765 -31.795 ;
        RECT 743.075 -32.125 743.405 -31.795 ;
        RECT 741.715 -32.125 742.045 -31.795 ;
        RECT 738.995 -32.125 739.325 -31.795 ;
        RECT 736.275 -32.125 736.605 -31.795 ;
        RECT 733.555 -32.125 733.885 -31.795 ;
        RECT 732.195 -32.125 732.525 -31.795 ;
        RECT 730.835 -32.125 731.165 -31.795 ;
        RECT 729.475 -32.125 729.805 -31.795 ;
        RECT 728.115 -32.125 728.445 -31.795 ;
        RECT 726.755 -32.125 727.085 -31.795 ;
        RECT 724.035 -32.125 724.365 -31.795 ;
        RECT 721.315 -32.125 721.645 -31.795 ;
        RECT 718.595 -32.125 718.925 -31.795 ;
        RECT 717.235 -32.125 717.565 -31.795 ;
        RECT 715.875 -32.125 716.205 -31.795 ;
        RECT 714.515 -32.125 714.845 -31.795 ;
        RECT 713.155 -32.125 713.485 -31.795 ;
        RECT 711.795 -32.125 712.125 -31.795 ;
        RECT 709.075 -32.125 709.405 -31.795 ;
        RECT 706.355 -32.125 706.685 -31.795 ;
        RECT 703.635 -32.125 703.965 -31.795 ;
        RECT 702.275 -32.125 702.605 -31.795 ;
        RECT 700.915 -32.125 701.245 -31.795 ;
        RECT 699.555 -32.125 699.885 -31.795 ;
        RECT 698.195 -32.125 698.525 -31.795 ;
        RECT 696.835 -32.125 697.165 -31.795 ;
        RECT 694.115 -32.125 694.445 -31.795 ;
        RECT 691.395 -32.125 691.725 -31.795 ;
        RECT 688.675 -32.125 689.005 -31.795 ;
        RECT 687.315 -32.125 687.645 -31.795 ;
        RECT 685.955 -32.125 686.285 -31.795 ;
        RECT 684.595 -32.125 684.925 -31.795 ;
        RECT 683.235 -32.125 683.565 -31.795 ;
        RECT 681.875 -32.125 682.205 -31.795 ;
        RECT 679.155 -32.125 679.485 -31.795 ;
        RECT 676.435 -32.125 676.765 -31.795 ;
        RECT 673.715 -32.125 674.045 -31.795 ;
        RECT 672.355 -32.125 672.685 -31.795 ;
        RECT 670.995 -32.125 671.325 -31.795 ;
        RECT 669.635 -32.125 669.965 -31.795 ;
        RECT 668.275 -32.125 668.605 -31.795 ;
        RECT 664.195 -32.125 664.525 -31.795 ;
        RECT 661.475 -32.125 661.805 -31.795 ;
        RECT 658.755 -32.125 659.085 -31.795 ;
        RECT 657.395 -32.125 657.725 -31.795 ;
        RECT 656.035 -32.125 656.365 -31.795 ;
        RECT 654.675 -32.125 655.005 -31.795 ;
        RECT 653.315 -32.125 653.645 -31.795 ;
        RECT 649.235 -32.125 649.565 -31.795 ;
        RECT 646.515 -32.125 646.845 -31.795 ;
        RECT 643.795 -32.125 644.125 -31.795 ;
        RECT 642.435 -32.125 642.765 -31.795 ;
        RECT 641.075 -32.125 641.405 -31.795 ;
        RECT 639.715 -32.125 640.045 -31.795 ;
        RECT 638.355 -32.125 638.685 -31.795 ;
        RECT 634.275 -32.125 634.605 -31.795 ;
        RECT 631.555 -32.125 631.885 -31.795 ;
        RECT 628.835 -32.125 629.165 -31.795 ;
        RECT 627.475 -32.125 627.805 -31.795 ;
        RECT 626.115 -32.125 626.445 -31.795 ;
        RECT 624.755 -32.125 625.085 -31.795 ;
        RECT 623.395 -32.125 623.725 -31.795 ;
        RECT 619.315 -32.125 619.645 -31.795 ;
        RECT 616.595 -32.125 616.925 -31.795 ;
        RECT 613.875 -32.125 614.205 -31.795 ;
        RECT 612.515 -32.125 612.845 -31.795 ;
        RECT 611.155 -32.125 611.485 -31.795 ;
        RECT 609.795 -32.125 610.125 -31.795 ;
        RECT 608.435 -32.125 608.765 -31.795 ;
        RECT 604.355 -32.125 604.685 -31.795 ;
        RECT 600.275 -32.125 600.605 -31.795 ;
        RECT 598.915 -32.125 599.245 -31.795 ;
        RECT 597.555 -32.125 597.885 -31.795 ;
        RECT 596.195 -32.125 596.525 -31.795 ;
        RECT 594.835 -32.125 595.165 -31.795 ;
        RECT 593.475 -32.125 593.805 -31.795 ;
        RECT 589.395 -32.125 589.725 -31.795 ;
        RECT 585.315 -32.125 585.645 -31.795 ;
        RECT 583.955 -32.125 584.285 -31.795 ;
        RECT 582.595 -32.125 582.925 -31.795 ;
        RECT 581.235 -32.125 581.565 -31.795 ;
        RECT 579.875 -32.125 580.205 -31.795 ;
        RECT 578.515 -32.125 578.845 -31.795 ;
        RECT 574.435 -32.125 574.765 -31.795 ;
        RECT 570.355 -32.125 570.685 -31.795 ;
        RECT 568.995 -32.125 569.325 -31.795 ;
        RECT 567.635 -32.125 567.965 -31.795 ;
        RECT 566.275 -32.125 566.605 -31.795 ;
        RECT 564.915 -32.125 565.245 -31.795 ;
        RECT 563.555 -32.125 563.885 -31.795 ;
        RECT 558.115 -32.125 558.445 -31.795 ;
        RECT 555.395 -32.125 555.725 -31.795 ;
        RECT 554.035 -32.125 554.365 -31.795 ;
        RECT 552.675 -32.125 553.005 -31.795 ;
        RECT 551.315 -32.125 551.645 -31.795 ;
        RECT 549.955 -32.125 550.285 -31.795 ;
        RECT 548.595 -32.125 548.925 -31.795 ;
        RECT 543.155 -32.125 543.485 -31.795 ;
        RECT 540.435 -32.125 540.765 -31.795 ;
        RECT 539.075 -32.125 539.405 -31.795 ;
        RECT 537.715 -32.125 538.045 -31.795 ;
        RECT 536.355 -32.125 536.685 -31.795 ;
        RECT 534.995 -32.125 535.325 -31.795 ;
        RECT 533.635 -32.125 533.965 -31.795 ;
        RECT 528.195 -32.125 528.525 -31.795 ;
        RECT 525.475 -32.125 525.805 -31.795 ;
        RECT 524.115 -32.125 524.445 -31.795 ;
        RECT 522.755 -32.125 523.085 -31.795 ;
        RECT 521.395 -32.125 521.725 -31.795 ;
        RECT 520.035 -32.125 520.365 -31.795 ;
        RECT 518.675 -32.125 519.005 -31.795 ;
        RECT 515.955 -32.125 516.285 -31.795 ;
        RECT 513.235 -32.125 513.565 -31.795 ;
        RECT 510.515 -32.125 510.845 -31.795 ;
        RECT 509.155 -32.125 509.485 -31.795 ;
        RECT 507.795 -32.125 508.125 -31.795 ;
        RECT 506.435 -32.125 506.765 -31.795 ;
        RECT 505.075 -32.125 505.405 -31.795 ;
        RECT 503.715 -32.125 504.045 -31.795 ;
        RECT 500.995 -32.125 501.325 -31.795 ;
        RECT 498.275 -32.125 498.605 -31.795 ;
        RECT 495.555 -32.125 495.885 -31.795 ;
        RECT 494.195 -32.125 494.525 -31.795 ;
        RECT 492.835 -32.125 493.165 -31.795 ;
        RECT 491.475 -32.125 491.805 -31.795 ;
        RECT 490.115 -32.125 490.445 -31.795 ;
        RECT 488.755 -32.125 489.085 -31.795 ;
        RECT 486.035 -32.125 486.365 -31.795 ;
        RECT 483.315 -32.125 483.645 -31.795 ;
        RECT 480.595 -32.125 480.925 -31.795 ;
        RECT 479.235 -32.125 479.565 -31.795 ;
        RECT 477.875 -32.125 478.205 -31.795 ;
        RECT 476.515 -32.125 476.845 -31.795 ;
        RECT 475.155 -32.125 475.485 -31.795 ;
        RECT 473.795 -32.125 474.125 -31.795 ;
        RECT 471.075 -32.125 471.405 -31.795 ;
        RECT 468.355 -32.125 468.685 -31.795 ;
        RECT 465.635 -32.125 465.965 -31.795 ;
        RECT 464.275 -32.125 464.605 -31.795 ;
        RECT 462.915 -32.125 463.245 -31.795 ;
        RECT 461.555 -32.125 461.885 -31.795 ;
        RECT 460.195 -32.125 460.525 -31.795 ;
        RECT 458.835 -32.125 459.165 -31.795 ;
        RECT 456.115 -32.125 456.445 -31.795 ;
        RECT 453.395 -32.125 453.725 -31.795 ;
        RECT 450.675 -32.125 451.005 -31.795 ;
        RECT 449.315 -32.125 449.645 -31.795 ;
        RECT 447.955 -32.125 448.285 -31.795 ;
        RECT 446.595 -32.125 446.925 -31.795 ;
        RECT 445.235 -32.125 445.565 -31.795 ;
        RECT 443.875 -32.125 444.205 -31.795 ;
        RECT 441.155 -32.125 441.485 -31.795 ;
        RECT 438.435 -32.125 438.765 -31.795 ;
        RECT 435.715 -32.125 436.045 -31.795 ;
        RECT 434.355 -32.125 434.685 -31.795 ;
        RECT 432.995 -32.125 433.325 -31.795 ;
        RECT 431.635 -32.125 431.965 -31.795 ;
        RECT 430.275 -32.125 430.605 -31.795 ;
        RECT 428.915 -32.125 429.245 -31.795 ;
        RECT 426.195 -32.125 426.525 -31.795 ;
        RECT 423.475 -32.125 423.805 -31.795 ;
        RECT 420.755 -32.125 421.085 -31.795 ;
        RECT 419.395 -32.125 419.725 -31.795 ;
        RECT 418.035 -32.125 418.365 -31.795 ;
        RECT 416.675 -32.125 417.005 -31.795 ;
        RECT 415.315 -32.125 415.645 -31.795 ;
        RECT 413.955 -32.125 414.285 -31.795 ;
        RECT 411.235 -32.125 411.565 -31.795 ;
        RECT 408.515 -32.125 408.845 -31.795 ;
        RECT 405.795 -32.125 406.125 -31.795 ;
        RECT 404.435 -32.125 404.765 -31.795 ;
        RECT 403.075 -32.125 403.405 -31.795 ;
        RECT 401.715 -32.125 402.045 -31.795 ;
        RECT 400.355 -32.125 400.685 -31.795 ;
        RECT 398.995 -32.125 399.325 -31.795 ;
        RECT 396.275 -32.125 396.605 -31.795 ;
        RECT 393.555 -32.125 393.885 -31.795 ;
        RECT 390.835 -32.125 391.165 -31.795 ;
        RECT 389.475 -32.125 389.805 -31.795 ;
        RECT 388.115 -32.125 388.445 -31.795 ;
        RECT 386.755 -32.125 387.085 -31.795 ;
        RECT 385.395 -32.125 385.725 -31.795 ;
        RECT 384.035 -32.125 384.365 -31.795 ;
        RECT 381.315 -32.125 381.645 -31.795 ;
        RECT 378.595 -32.125 378.925 -31.795 ;
        RECT 375.875 -32.125 376.205 -31.795 ;
        RECT 374.515 -32.125 374.845 -31.795 ;
        RECT 373.155 -32.125 373.485 -31.795 ;
        RECT 371.795 -32.125 372.125 -31.795 ;
        RECT 370.435 -32.125 370.765 -31.795 ;
        RECT 369.075 -32.125 369.405 -31.795 ;
        RECT 366.355 -32.125 366.685 -31.795 ;
        RECT 363.635 -32.125 363.965 -31.795 ;
        RECT 360.915 -32.125 361.245 -31.795 ;
        RECT 359.555 -32.125 359.885 -31.795 ;
        RECT 358.195 -32.125 358.525 -31.795 ;
        RECT 356.835 -32.125 357.165 -31.795 ;
        RECT 355.475 -32.125 355.805 -31.795 ;
        RECT 354.115 -32.125 354.445 -31.795 ;
        RECT 351.395 -32.125 351.725 -31.795 ;
        RECT 348.675 -32.125 349.005 -31.795 ;
        RECT 345.955 -32.125 346.285 -31.795 ;
        RECT 344.595 -32.125 344.925 -31.795 ;
        RECT 343.235 -32.125 343.565 -31.795 ;
        RECT 341.875 -32.125 342.205 -31.795 ;
        RECT 340.515 -32.125 340.845 -31.795 ;
        RECT 339.155 -32.125 339.485 -31.795 ;
        RECT 336.435 -32.125 336.765 -31.795 ;
        RECT 333.715 -32.125 334.045 -31.795 ;
        RECT 330.995 -32.125 331.325 -31.795 ;
        RECT 329.635 -32.125 329.965 -31.795 ;
        RECT 328.275 -32.125 328.605 -31.795 ;
        RECT 326.915 -32.125 327.245 -31.795 ;
        RECT 325.555 -32.125 325.885 -31.795 ;
        RECT 321.475 -32.125 321.805 -31.795 ;
        RECT 318.755 -32.125 319.085 -31.795 ;
        RECT 316.035 -32.125 316.365 -31.795 ;
        RECT 314.675 -32.125 315.005 -31.795 ;
        RECT 313.315 -32.125 313.645 -31.795 ;
        RECT 311.955 -32.125 312.285 -31.795 ;
        RECT 310.595 -32.125 310.925 -31.795 ;
        RECT 306.515 -32.125 306.845 -31.795 ;
        RECT 303.795 -32.125 304.125 -31.795 ;
        RECT 301.075 -32.125 301.405 -31.795 ;
        RECT 299.715 -32.125 300.045 -31.795 ;
        RECT 298.355 -32.125 298.685 -31.795 ;
        RECT 296.995 -32.125 297.325 -31.795 ;
        RECT 295.635 -32.125 295.965 -31.795 ;
        RECT 291.555 -32.125 291.885 -31.795 ;
        RECT 288.835 -32.125 289.165 -31.795 ;
        RECT 286.115 -32.125 286.445 -31.795 ;
        RECT 284.755 -32.125 285.085 -31.795 ;
        RECT 283.395 -32.125 283.725 -31.795 ;
        RECT 282.035 -32.125 282.365 -31.795 ;
        RECT 280.675 -32.125 281.005 -31.795 ;
        RECT 276.595 -32.125 276.925 -31.795 ;
        RECT 273.875 -32.125 274.205 -31.795 ;
        RECT 272.515 -32.125 272.845 -31.795 ;
        RECT 271.155 -32.125 271.485 -31.795 ;
        RECT 269.795 -32.125 270.125 -31.795 ;
        RECT 268.435 -32.125 268.765 -31.795 ;
        RECT 267.075 -32.125 267.405 -31.795 ;
        RECT 265.715 -32.125 266.045 -31.795 ;
        RECT 261.635 -32.125 261.965 -31.795 ;
        RECT 257.555 -32.125 257.885 -31.795 ;
        RECT 256.195 -32.125 256.525 -31.795 ;
        RECT 254.835 -32.125 255.165 -31.795 ;
        RECT 253.475 -32.125 253.805 -31.795 ;
        RECT 252.115 -32.125 252.445 -31.795 ;
        RECT 250.755 -32.125 251.085 -31.795 ;
        RECT 246.675 -32.125 247.005 -31.795 ;
        RECT 242.595 -32.125 242.925 -31.795 ;
        RECT 241.235 -32.125 241.565 -31.795 ;
        RECT 239.875 -32.125 240.205 -31.795 ;
        RECT 238.515 -32.125 238.845 -31.795 ;
        RECT 237.155 -32.125 237.485 -31.795 ;
        RECT 235.795 -32.125 236.125 -31.795 ;
        RECT 231.715 -32.125 232.045 -31.795 ;
        RECT 227.635 -32.125 227.965 -31.795 ;
        RECT 226.275 -32.125 226.605 -31.795 ;
        RECT 224.915 -32.125 225.245 -31.795 ;
        RECT 223.555 -32.125 223.885 -31.795 ;
        RECT 222.195 -32.125 222.525 -31.795 ;
        RECT 220.835 -32.125 221.165 -31.795 ;
        RECT 215.395 -32.125 215.725 -31.795 ;
        RECT 212.675 -32.125 213.005 -31.795 ;
        RECT 211.315 -32.125 211.645 -31.795 ;
        RECT 209.955 -32.125 210.285 -31.795 ;
        RECT 208.595 -32.125 208.925 -31.795 ;
        RECT 207.235 -32.125 207.565 -31.795 ;
        RECT 205.875 -32.125 206.205 -31.795 ;
        RECT 200.435 -32.125 200.765 -31.795 ;
        RECT 197.715 -32.125 198.045 -31.795 ;
        RECT 196.355 -32.125 196.685 -31.795 ;
        RECT 194.995 -32.125 195.325 -31.795 ;
        RECT 193.635 -32.125 193.965 -31.795 ;
        RECT 192.275 -32.125 192.605 -31.795 ;
        RECT 190.915 -32.125 191.245 -31.795 ;
        RECT 185.475 -32.125 185.805 -31.795 ;
        RECT 182.755 -32.125 183.085 -31.795 ;
        RECT 181.395 -32.125 181.725 -31.795 ;
        RECT 180.035 -32.125 180.365 -31.795 ;
        RECT 178.675 -32.125 179.005 -31.795 ;
        RECT 177.315 -32.125 177.645 -31.795 ;
        RECT 175.955 -32.125 176.285 -31.795 ;
        RECT 173.235 -32.125 173.565 -31.795 ;
        RECT 170.515 -32.125 170.845 -31.795 ;
        RECT 167.795 -32.125 168.125 -31.795 ;
        RECT 166.435 -32.125 166.765 -31.795 ;
        RECT 165.075 -32.125 165.405 -31.795 ;
        RECT 163.715 -32.125 164.045 -31.795 ;
        RECT 162.355 -32.125 162.685 -31.795 ;
        RECT 160.995 -32.125 161.325 -31.795 ;
        RECT 158.275 -32.125 158.605 -31.795 ;
        RECT 155.555 -32.125 155.885 -31.795 ;
        RECT 152.835 -32.125 153.165 -31.795 ;
        RECT 151.475 -32.125 151.805 -31.795 ;
        RECT 150.115 -32.125 150.445 -31.795 ;
        RECT 148.755 -32.125 149.085 -31.795 ;
        RECT 147.395 -32.125 147.725 -31.795 ;
        RECT 146.035 -32.125 146.365 -31.795 ;
        RECT 143.315 -32.125 143.645 -31.795 ;
        RECT 140.595 -32.125 140.925 -31.795 ;
        RECT 137.875 -32.125 138.205 -31.795 ;
        RECT 136.515 -32.125 136.845 -31.795 ;
        RECT 135.155 -32.125 135.485 -31.795 ;
        RECT 133.795 -32.125 134.125 -31.795 ;
        RECT 132.435 -32.125 132.765 -31.795 ;
        RECT 131.075 -32.125 131.405 -31.795 ;
        RECT 128.355 -32.125 128.685 -31.795 ;
        RECT 125.635 -32.125 125.965 -31.795 ;
        RECT 122.915 -32.125 123.245 -31.795 ;
        RECT 121.555 -32.125 121.885 -31.795 ;
        RECT 120.195 -32.125 120.525 -31.795 ;
        RECT 118.835 -32.125 119.165 -31.795 ;
        RECT 117.475 -32.125 117.805 -31.795 ;
        RECT 116.115 -32.125 116.445 -31.795 ;
        RECT 113.395 -32.125 113.725 -31.795 ;
        RECT 110.675 -32.125 111.005 -31.795 ;
        RECT 107.955 -32.125 108.285 -31.795 ;
        RECT 106.595 -32.125 106.925 -31.795 ;
        RECT 105.235 -32.125 105.565 -31.795 ;
        RECT 103.875 -32.125 104.205 -31.795 ;
        RECT 102.515 -32.125 102.845 -31.795 ;
        RECT 101.155 -32.125 101.485 -31.795 ;
        RECT 98.435 -32.125 98.765 -31.795 ;
        RECT 95.715 -32.125 96.045 -31.795 ;
        RECT 92.995 -32.125 93.325 -31.795 ;
        RECT 91.635 -32.125 91.965 -31.795 ;
        RECT 90.275 -32.125 90.605 -31.795 ;
        RECT 88.915 -32.125 89.245 -31.795 ;
        RECT 87.555 -32.125 87.885 -31.795 ;
        RECT 86.195 -32.125 86.525 -31.795 ;
        RECT 83.475 -32.125 83.805 -31.795 ;
        RECT 80.755 -32.125 81.085 -31.795 ;
        RECT 78.035 -32.125 78.365 -31.795 ;
        RECT 76.675 -32.125 77.005 -31.795 ;
        RECT 75.315 -32.125 75.645 -31.795 ;
        RECT 73.955 -32.125 74.285 -31.795 ;
        RECT 72.595 -32.125 72.925 -31.795 ;
        RECT 71.235 -32.125 71.565 -31.795 ;
        RECT 68.515 -32.125 68.845 -31.795 ;
        RECT 65.795 -32.125 66.125 -31.795 ;
        RECT 63.075 -32.125 63.405 -31.795 ;
        RECT 61.715 -32.125 62.045 -31.795 ;
        RECT 60.355 -32.125 60.685 -31.795 ;
        RECT 58.995 -32.125 59.325 -31.795 ;
        RECT 57.635 -32.125 57.965 -31.795 ;
        RECT 56.275 -32.125 56.605 -31.795 ;
        RECT 53.555 -32.125 53.885 -31.795 ;
        RECT 50.835 -32.125 51.165 -31.795 ;
        RECT 48.115 -32.125 48.445 -31.795 ;
        RECT 46.755 -32.125 47.085 -31.795 ;
        RECT 45.395 -32.125 45.725 -31.795 ;
        RECT 44.035 -32.125 44.365 -31.795 ;
        RECT 42.675 -32.125 43.005 -31.795 ;
        RECT 41.315 -32.125 41.645 -31.795 ;
        RECT 38.595 -32.125 38.925 -31.795 ;
        RECT 35.875 -32.125 36.205 -31.795 ;
        RECT 33.155 -32.125 33.485 -31.795 ;
        RECT 31.795 -32.125 32.125 -31.795 ;
        RECT 30.435 -32.125 30.765 -31.795 ;
        RECT 29.075 -32.125 29.405 -31.795 ;
        RECT 27.715 -32.125 28.045 -31.795 ;
        RECT 26.355 -32.125 26.685 -31.795 ;
        RECT 23.635 -32.125 23.965 -31.795 ;
        RECT 20.915 -32.125 21.245 -31.795 ;
        RECT 18.195 -32.125 18.525 -31.795 ;
        RECT 16.835 -32.125 17.165 -31.795 ;
        RECT 15.475 -32.125 15.805 -31.795 ;
        RECT 14.115 -32.125 14.445 -31.795 ;
        RECT 12.755 -32.125 13.085 -31.795 ;
        RECT 11.395 -32.125 11.725 -31.795 ;
        RECT 8.675 -32.125 9.005 -31.795 ;
        RECT 7.315 -32.125 7.645 -31.795 ;
        RECT 5.955 -32.125 6.285 -31.795 ;
        RECT 4.595 -32.125 4.925 -31.795 ;
        RECT 3.235 -32.125 3.565 -31.795 ;
        RECT 1.875 -32.125 2.205 -31.795 ;
        RECT 0.515 -32.125 0.845 -31.795 ;
        RECT -0.845 -32.125 -0.515 -31.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -33.48 954.88 -33.16 ;
        RECT 953.875 -33.485 954.205 -33.155 ;
        RECT 952.515 -33.485 952.845 -33.155 ;
        RECT 951.155 -33.485 951.485 -33.155 ;
        RECT 949.795 -33.485 950.125 -33.155 ;
        RECT 947.075 -33.485 947.405 -33.155 ;
        RECT 945.715 -33.485 946.045 -33.155 ;
        RECT 944.355 -33.485 944.685 -33.155 ;
        RECT 942.995 -33.485 943.325 -33.155 ;
        RECT 941.635 -33.485 941.965 -33.155 ;
        RECT 940.275 -33.485 940.605 -33.155 ;
        RECT 938.915 -33.485 939.245 -33.155 ;
        RECT 937.555 -33.485 937.885 -33.155 ;
        RECT 936.195 -33.485 936.525 -33.155 ;
        RECT 932.115 -33.485 932.445 -33.155 ;
        RECT 928.035 -33.485 928.365 -33.155 ;
        RECT 926.675 -33.485 927.005 -33.155 ;
        RECT 925.315 -33.485 925.645 -33.155 ;
        RECT 923.955 -33.485 924.285 -33.155 ;
        RECT 922.595 -33.485 922.925 -33.155 ;
        RECT 921.235 -33.485 921.565 -33.155 ;
        RECT 917.155 -33.485 917.485 -33.155 ;
        RECT 913.075 -33.485 913.405 -33.155 ;
        RECT 911.715 -33.485 912.045 -33.155 ;
        RECT 910.355 -33.485 910.685 -33.155 ;
        RECT 908.995 -33.485 909.325 -33.155 ;
        RECT 907.635 -33.485 907.965 -33.155 ;
        RECT 906.275 -33.485 906.605 -33.155 ;
        RECT 902.195 -33.485 902.525 -33.155 ;
        RECT 900.835 -33.485 901.165 -33.155 ;
        RECT 898.115 -33.485 898.445 -33.155 ;
        RECT 896.755 -33.485 897.085 -33.155 ;
        RECT 895.395 -33.485 895.725 -33.155 ;
        RECT 894.035 -33.485 894.365 -33.155 ;
        RECT 892.675 -33.485 893.005 -33.155 ;
        RECT 891.315 -33.485 891.645 -33.155 ;
        RECT 885.875 -33.485 886.205 -33.155 ;
        RECT 883.155 -33.485 883.485 -33.155 ;
        RECT 881.795 -33.485 882.125 -33.155 ;
        RECT 880.435 -33.485 880.765 -33.155 ;
        RECT 879.075 -33.485 879.405 -33.155 ;
        RECT 877.715 -33.485 878.045 -33.155 ;
        RECT 876.355 -33.485 876.685 -33.155 ;
        RECT 870.915 -33.485 871.245 -33.155 ;
        RECT 868.195 -33.485 868.525 -33.155 ;
        RECT 866.835 -33.485 867.165 -33.155 ;
        RECT 865.475 -33.485 865.805 -33.155 ;
        RECT 864.115 -33.485 864.445 -33.155 ;
        RECT 862.755 -33.485 863.085 -33.155 ;
        RECT 861.395 -33.485 861.725 -33.155 ;
        RECT 855.955 -33.485 856.285 -33.155 ;
        RECT 853.235 -33.485 853.565 -33.155 ;
        RECT 851.875 -33.485 852.205 -33.155 ;
        RECT 850.515 -33.485 850.845 -33.155 ;
        RECT 849.155 -33.485 849.485 -33.155 ;
        RECT 847.795 -33.485 848.125 -33.155 ;
        RECT 846.435 -33.485 846.765 -33.155 ;
        RECT 843.715 -33.485 844.045 -33.155 ;
        RECT 840.995 -33.485 841.325 -33.155 ;
        RECT 838.275 -33.485 838.605 -33.155 ;
        RECT 836.915 -33.485 837.245 -33.155 ;
        RECT 835.555 -33.485 835.885 -33.155 ;
        RECT 834.195 -33.485 834.525 -33.155 ;
        RECT 832.835 -33.485 833.165 -33.155 ;
        RECT 831.475 -33.485 831.805 -33.155 ;
        RECT 828.755 -33.485 829.085 -33.155 ;
        RECT 826.035 -33.485 826.365 -33.155 ;
        RECT 823.315 -33.485 823.645 -33.155 ;
        RECT 821.955 -33.485 822.285 -33.155 ;
        RECT 820.595 -33.485 820.925 -33.155 ;
        RECT 819.235 -33.485 819.565 -33.155 ;
        RECT 817.875 -33.485 818.205 -33.155 ;
        RECT 816.515 -33.485 816.845 -33.155 ;
        RECT 813.795 -33.485 814.125 -33.155 ;
        RECT 811.075 -33.485 811.405 -33.155 ;
        RECT 808.355 -33.485 808.685 -33.155 ;
        RECT 806.995 -33.485 807.325 -33.155 ;
        RECT 805.635 -33.485 805.965 -33.155 ;
        RECT 804.275 -33.485 804.605 -33.155 ;
        RECT 802.915 -33.485 803.245 -33.155 ;
        RECT 801.555 -33.485 801.885 -33.155 ;
        RECT 798.835 -33.485 799.165 -33.155 ;
        RECT 796.115 -33.485 796.445 -33.155 ;
        RECT 793.395 -33.485 793.725 -33.155 ;
        RECT 792.035 -33.485 792.365 -33.155 ;
        RECT 790.675 -33.485 791.005 -33.155 ;
        RECT 789.315 -33.485 789.645 -33.155 ;
        RECT 787.955 -33.485 788.285 -33.155 ;
        RECT 786.595 -33.485 786.925 -33.155 ;
        RECT 783.875 -33.485 784.205 -33.155 ;
        RECT 781.155 -33.485 781.485 -33.155 ;
        RECT 778.435 -33.485 778.765 -33.155 ;
        RECT 777.075 -33.485 777.405 -33.155 ;
        RECT 775.715 -33.485 776.045 -33.155 ;
        RECT 774.355 -33.485 774.685 -33.155 ;
        RECT 772.995 -33.485 773.325 -33.155 ;
        RECT 771.635 -33.485 771.965 -33.155 ;
        RECT 768.915 -33.485 769.245 -33.155 ;
        RECT 766.195 -33.485 766.525 -33.155 ;
        RECT 763.475 -33.485 763.805 -33.155 ;
        RECT 762.115 -33.485 762.445 -33.155 ;
        RECT 760.755 -33.485 761.085 -33.155 ;
        RECT 759.395 -33.485 759.725 -33.155 ;
        RECT 758.035 -33.485 758.365 -33.155 ;
        RECT 756.675 -33.485 757.005 -33.155 ;
        RECT 753.955 -33.485 754.285 -33.155 ;
        RECT 751.235 -33.485 751.565 -33.155 ;
        RECT 748.515 -33.485 748.845 -33.155 ;
        RECT 747.155 -33.485 747.485 -33.155 ;
        RECT 745.795 -33.485 746.125 -33.155 ;
        RECT 744.435 -33.485 744.765 -33.155 ;
        RECT 743.075 -33.485 743.405 -33.155 ;
        RECT 741.715 -33.485 742.045 -33.155 ;
        RECT 738.995 -33.485 739.325 -33.155 ;
        RECT 736.275 -33.485 736.605 -33.155 ;
        RECT 733.555 -33.485 733.885 -33.155 ;
        RECT 732.195 -33.485 732.525 -33.155 ;
        RECT 730.835 -33.485 731.165 -33.155 ;
        RECT 729.475 -33.485 729.805 -33.155 ;
        RECT 728.115 -33.485 728.445 -33.155 ;
        RECT 726.755 -33.485 727.085 -33.155 ;
        RECT 724.035 -33.485 724.365 -33.155 ;
        RECT 721.315 -33.485 721.645 -33.155 ;
        RECT 718.595 -33.485 718.925 -33.155 ;
        RECT 717.235 -33.485 717.565 -33.155 ;
        RECT 715.875 -33.485 716.205 -33.155 ;
        RECT 714.515 -33.485 714.845 -33.155 ;
        RECT 713.155 -33.485 713.485 -33.155 ;
        RECT 711.795 -33.485 712.125 -33.155 ;
        RECT 709.075 -33.485 709.405 -33.155 ;
        RECT 706.355 -33.485 706.685 -33.155 ;
        RECT 703.635 -33.485 703.965 -33.155 ;
        RECT 702.275 -33.485 702.605 -33.155 ;
        RECT 700.915 -33.485 701.245 -33.155 ;
        RECT 699.555 -33.485 699.885 -33.155 ;
        RECT 698.195 -33.485 698.525 -33.155 ;
        RECT 696.835 -33.485 697.165 -33.155 ;
        RECT 694.115 -33.485 694.445 -33.155 ;
        RECT 691.395 -33.485 691.725 -33.155 ;
        RECT 688.675 -33.485 689.005 -33.155 ;
        RECT 687.315 -33.485 687.645 -33.155 ;
        RECT 685.955 -33.485 686.285 -33.155 ;
        RECT 684.595 -33.485 684.925 -33.155 ;
        RECT 683.235 -33.485 683.565 -33.155 ;
        RECT 681.875 -33.485 682.205 -33.155 ;
        RECT 679.155 -33.485 679.485 -33.155 ;
        RECT 676.435 -33.485 676.765 -33.155 ;
        RECT 673.715 -33.485 674.045 -33.155 ;
        RECT 672.355 -33.485 672.685 -33.155 ;
        RECT 670.995 -33.485 671.325 -33.155 ;
        RECT 669.635 -33.485 669.965 -33.155 ;
        RECT 668.275 -33.485 668.605 -33.155 ;
        RECT 664.195 -33.485 664.525 -33.155 ;
        RECT 661.475 -33.485 661.805 -33.155 ;
        RECT 658.755 -33.485 659.085 -33.155 ;
        RECT 657.395 -33.485 657.725 -33.155 ;
        RECT 656.035 -33.485 656.365 -33.155 ;
        RECT 654.675 -33.485 655.005 -33.155 ;
        RECT 653.315 -33.485 653.645 -33.155 ;
        RECT 649.235 -33.485 649.565 -33.155 ;
        RECT 646.515 -33.485 646.845 -33.155 ;
        RECT 643.795 -33.485 644.125 -33.155 ;
        RECT 642.435 -33.485 642.765 -33.155 ;
        RECT 641.075 -33.485 641.405 -33.155 ;
        RECT 639.715 -33.485 640.045 -33.155 ;
        RECT 638.355 -33.485 638.685 -33.155 ;
        RECT 634.275 -33.485 634.605 -33.155 ;
        RECT 631.555 -33.485 631.885 -33.155 ;
        RECT 628.835 -33.485 629.165 -33.155 ;
        RECT 627.475 -33.485 627.805 -33.155 ;
        RECT 626.115 -33.485 626.445 -33.155 ;
        RECT 624.755 -33.485 625.085 -33.155 ;
        RECT 623.395 -33.485 623.725 -33.155 ;
        RECT 619.315 -33.485 619.645 -33.155 ;
        RECT 616.595 -33.485 616.925 -33.155 ;
        RECT 613.875 -33.485 614.205 -33.155 ;
        RECT 612.515 -33.485 612.845 -33.155 ;
        RECT 611.155 -33.485 611.485 -33.155 ;
        RECT 609.795 -33.485 610.125 -33.155 ;
        RECT 608.435 -33.485 608.765 -33.155 ;
        RECT 604.355 -33.485 604.685 -33.155 ;
        RECT 600.275 -33.485 600.605 -33.155 ;
        RECT 598.915 -33.485 599.245 -33.155 ;
        RECT 597.555 -33.485 597.885 -33.155 ;
        RECT 596.195 -33.485 596.525 -33.155 ;
        RECT 594.835 -33.485 595.165 -33.155 ;
        RECT 593.475 -33.485 593.805 -33.155 ;
        RECT 589.395 -33.485 589.725 -33.155 ;
        RECT 585.315 -33.485 585.645 -33.155 ;
        RECT 583.955 -33.485 584.285 -33.155 ;
        RECT 582.595 -33.485 582.925 -33.155 ;
        RECT 581.235 -33.485 581.565 -33.155 ;
        RECT 579.875 -33.485 580.205 -33.155 ;
        RECT 578.515 -33.485 578.845 -33.155 ;
        RECT 574.435 -33.485 574.765 -33.155 ;
        RECT 570.355 -33.485 570.685 -33.155 ;
        RECT 568.995 -33.485 569.325 -33.155 ;
        RECT 567.635 -33.485 567.965 -33.155 ;
        RECT 566.275 -33.485 566.605 -33.155 ;
        RECT 564.915 -33.485 565.245 -33.155 ;
        RECT 563.555 -33.485 563.885 -33.155 ;
        RECT 558.115 -33.485 558.445 -33.155 ;
        RECT 555.395 -33.485 555.725 -33.155 ;
        RECT 554.035 -33.485 554.365 -33.155 ;
        RECT 552.675 -33.485 553.005 -33.155 ;
        RECT 551.315 -33.485 551.645 -33.155 ;
        RECT 549.955 -33.485 550.285 -33.155 ;
        RECT 548.595 -33.485 548.925 -33.155 ;
        RECT 543.155 -33.485 543.485 -33.155 ;
        RECT 540.435 -33.485 540.765 -33.155 ;
        RECT 539.075 -33.485 539.405 -33.155 ;
        RECT 537.715 -33.485 538.045 -33.155 ;
        RECT 536.355 -33.485 536.685 -33.155 ;
        RECT 534.995 -33.485 535.325 -33.155 ;
        RECT 533.635 -33.485 533.965 -33.155 ;
        RECT 528.195 -33.485 528.525 -33.155 ;
        RECT 525.475 -33.485 525.805 -33.155 ;
        RECT 524.115 -33.485 524.445 -33.155 ;
        RECT 522.755 -33.485 523.085 -33.155 ;
        RECT 521.395 -33.485 521.725 -33.155 ;
        RECT 520.035 -33.485 520.365 -33.155 ;
        RECT 518.675 -33.485 519.005 -33.155 ;
        RECT 515.955 -33.485 516.285 -33.155 ;
        RECT 513.235 -33.485 513.565 -33.155 ;
        RECT 510.515 -33.485 510.845 -33.155 ;
        RECT 509.155 -33.485 509.485 -33.155 ;
        RECT 507.795 -33.485 508.125 -33.155 ;
        RECT 506.435 -33.485 506.765 -33.155 ;
        RECT 505.075 -33.485 505.405 -33.155 ;
        RECT 503.715 -33.485 504.045 -33.155 ;
        RECT 500.995 -33.485 501.325 -33.155 ;
        RECT 498.275 -33.485 498.605 -33.155 ;
        RECT 495.555 -33.485 495.885 -33.155 ;
        RECT 494.195 -33.485 494.525 -33.155 ;
        RECT 492.835 -33.485 493.165 -33.155 ;
        RECT 491.475 -33.485 491.805 -33.155 ;
        RECT 490.115 -33.485 490.445 -33.155 ;
        RECT 488.755 -33.485 489.085 -33.155 ;
        RECT 486.035 -33.485 486.365 -33.155 ;
        RECT 483.315 -33.485 483.645 -33.155 ;
        RECT 480.595 -33.485 480.925 -33.155 ;
        RECT 479.235 -33.485 479.565 -33.155 ;
        RECT 477.875 -33.485 478.205 -33.155 ;
        RECT 476.515 -33.485 476.845 -33.155 ;
        RECT 475.155 -33.485 475.485 -33.155 ;
        RECT 473.795 -33.485 474.125 -33.155 ;
        RECT 471.075 -33.485 471.405 -33.155 ;
        RECT 468.355 -33.485 468.685 -33.155 ;
        RECT 465.635 -33.485 465.965 -33.155 ;
        RECT 464.275 -33.485 464.605 -33.155 ;
        RECT 462.915 -33.485 463.245 -33.155 ;
        RECT 461.555 -33.485 461.885 -33.155 ;
        RECT 460.195 -33.485 460.525 -33.155 ;
        RECT 458.835 -33.485 459.165 -33.155 ;
        RECT 456.115 -33.485 456.445 -33.155 ;
        RECT 453.395 -33.485 453.725 -33.155 ;
        RECT 450.675 -33.485 451.005 -33.155 ;
        RECT 449.315 -33.485 449.645 -33.155 ;
        RECT 447.955 -33.485 448.285 -33.155 ;
        RECT 446.595 -33.485 446.925 -33.155 ;
        RECT 445.235 -33.485 445.565 -33.155 ;
        RECT 443.875 -33.485 444.205 -33.155 ;
        RECT 441.155 -33.485 441.485 -33.155 ;
        RECT 438.435 -33.485 438.765 -33.155 ;
        RECT 435.715 -33.485 436.045 -33.155 ;
        RECT 434.355 -33.485 434.685 -33.155 ;
        RECT 432.995 -33.485 433.325 -33.155 ;
        RECT 431.635 -33.485 431.965 -33.155 ;
        RECT 430.275 -33.485 430.605 -33.155 ;
        RECT 428.915 -33.485 429.245 -33.155 ;
        RECT 426.195 -33.485 426.525 -33.155 ;
        RECT 423.475 -33.485 423.805 -33.155 ;
        RECT 420.755 -33.485 421.085 -33.155 ;
        RECT 419.395 -33.485 419.725 -33.155 ;
        RECT 418.035 -33.485 418.365 -33.155 ;
        RECT 416.675 -33.485 417.005 -33.155 ;
        RECT 415.315 -33.485 415.645 -33.155 ;
        RECT 413.955 -33.485 414.285 -33.155 ;
        RECT 411.235 -33.485 411.565 -33.155 ;
        RECT 408.515 -33.485 408.845 -33.155 ;
        RECT 405.795 -33.485 406.125 -33.155 ;
        RECT 404.435 -33.485 404.765 -33.155 ;
        RECT 403.075 -33.485 403.405 -33.155 ;
        RECT 401.715 -33.485 402.045 -33.155 ;
        RECT 400.355 -33.485 400.685 -33.155 ;
        RECT 398.995 -33.485 399.325 -33.155 ;
        RECT 396.275 -33.485 396.605 -33.155 ;
        RECT 393.555 -33.485 393.885 -33.155 ;
        RECT 390.835 -33.485 391.165 -33.155 ;
        RECT 389.475 -33.485 389.805 -33.155 ;
        RECT 388.115 -33.485 388.445 -33.155 ;
        RECT 386.755 -33.485 387.085 -33.155 ;
        RECT 385.395 -33.485 385.725 -33.155 ;
        RECT 384.035 -33.485 384.365 -33.155 ;
        RECT 381.315 -33.485 381.645 -33.155 ;
        RECT 378.595 -33.485 378.925 -33.155 ;
        RECT 375.875 -33.485 376.205 -33.155 ;
        RECT 374.515 -33.485 374.845 -33.155 ;
        RECT 373.155 -33.485 373.485 -33.155 ;
        RECT 371.795 -33.485 372.125 -33.155 ;
        RECT 370.435 -33.485 370.765 -33.155 ;
        RECT 369.075 -33.485 369.405 -33.155 ;
        RECT 366.355 -33.485 366.685 -33.155 ;
        RECT 363.635 -33.485 363.965 -33.155 ;
        RECT 360.915 -33.485 361.245 -33.155 ;
        RECT 359.555 -33.485 359.885 -33.155 ;
        RECT 358.195 -33.485 358.525 -33.155 ;
        RECT 356.835 -33.485 357.165 -33.155 ;
        RECT 355.475 -33.485 355.805 -33.155 ;
        RECT 354.115 -33.485 354.445 -33.155 ;
        RECT 351.395 -33.485 351.725 -33.155 ;
        RECT 348.675 -33.485 349.005 -33.155 ;
        RECT 345.955 -33.485 346.285 -33.155 ;
        RECT 344.595 -33.485 344.925 -33.155 ;
        RECT 343.235 -33.485 343.565 -33.155 ;
        RECT 341.875 -33.485 342.205 -33.155 ;
        RECT 340.515 -33.485 340.845 -33.155 ;
        RECT 339.155 -33.485 339.485 -33.155 ;
        RECT 336.435 -33.485 336.765 -33.155 ;
        RECT 333.715 -33.485 334.045 -33.155 ;
        RECT 330.995 -33.485 331.325 -33.155 ;
        RECT 329.635 -33.485 329.965 -33.155 ;
        RECT 328.275 -33.485 328.605 -33.155 ;
        RECT 326.915 -33.485 327.245 -33.155 ;
        RECT 325.555 -33.485 325.885 -33.155 ;
        RECT 321.475 -33.485 321.805 -33.155 ;
        RECT 318.755 -33.485 319.085 -33.155 ;
        RECT 316.035 -33.485 316.365 -33.155 ;
        RECT 314.675 -33.485 315.005 -33.155 ;
        RECT 313.315 -33.485 313.645 -33.155 ;
        RECT 311.955 -33.485 312.285 -33.155 ;
        RECT 310.595 -33.485 310.925 -33.155 ;
        RECT 306.515 -33.485 306.845 -33.155 ;
        RECT 303.795 -33.485 304.125 -33.155 ;
        RECT 301.075 -33.485 301.405 -33.155 ;
        RECT 299.715 -33.485 300.045 -33.155 ;
        RECT 298.355 -33.485 298.685 -33.155 ;
        RECT 296.995 -33.485 297.325 -33.155 ;
        RECT 295.635 -33.485 295.965 -33.155 ;
        RECT 291.555 -33.485 291.885 -33.155 ;
        RECT 288.835 -33.485 289.165 -33.155 ;
        RECT 286.115 -33.485 286.445 -33.155 ;
        RECT 284.755 -33.485 285.085 -33.155 ;
        RECT 283.395 -33.485 283.725 -33.155 ;
        RECT 282.035 -33.485 282.365 -33.155 ;
        RECT 280.675 -33.485 281.005 -33.155 ;
        RECT 276.595 -33.485 276.925 -33.155 ;
        RECT 273.875 -33.485 274.205 -33.155 ;
        RECT 272.515 -33.485 272.845 -33.155 ;
        RECT 271.155 -33.485 271.485 -33.155 ;
        RECT 269.795 -33.485 270.125 -33.155 ;
        RECT 268.435 -33.485 268.765 -33.155 ;
        RECT 267.075 -33.485 267.405 -33.155 ;
        RECT 265.715 -33.485 266.045 -33.155 ;
        RECT 261.635 -33.485 261.965 -33.155 ;
        RECT 257.555 -33.485 257.885 -33.155 ;
        RECT 256.195 -33.485 256.525 -33.155 ;
        RECT 254.835 -33.485 255.165 -33.155 ;
        RECT 253.475 -33.485 253.805 -33.155 ;
        RECT 252.115 -33.485 252.445 -33.155 ;
        RECT 250.755 -33.485 251.085 -33.155 ;
        RECT 246.675 -33.485 247.005 -33.155 ;
        RECT 242.595 -33.485 242.925 -33.155 ;
        RECT 241.235 -33.485 241.565 -33.155 ;
        RECT 239.875 -33.485 240.205 -33.155 ;
        RECT 238.515 -33.485 238.845 -33.155 ;
        RECT 237.155 -33.485 237.485 -33.155 ;
        RECT 235.795 -33.485 236.125 -33.155 ;
        RECT 231.715 -33.485 232.045 -33.155 ;
        RECT 227.635 -33.485 227.965 -33.155 ;
        RECT 226.275 -33.485 226.605 -33.155 ;
        RECT 224.915 -33.485 225.245 -33.155 ;
        RECT 223.555 -33.485 223.885 -33.155 ;
        RECT 222.195 -33.485 222.525 -33.155 ;
        RECT 220.835 -33.485 221.165 -33.155 ;
        RECT 215.395 -33.485 215.725 -33.155 ;
        RECT 212.675 -33.485 213.005 -33.155 ;
        RECT 211.315 -33.485 211.645 -33.155 ;
        RECT 209.955 -33.485 210.285 -33.155 ;
        RECT 208.595 -33.485 208.925 -33.155 ;
        RECT 207.235 -33.485 207.565 -33.155 ;
        RECT 205.875 -33.485 206.205 -33.155 ;
        RECT 200.435 -33.485 200.765 -33.155 ;
        RECT 197.715 -33.485 198.045 -33.155 ;
        RECT 196.355 -33.485 196.685 -33.155 ;
        RECT 194.995 -33.485 195.325 -33.155 ;
        RECT 193.635 -33.485 193.965 -33.155 ;
        RECT 192.275 -33.485 192.605 -33.155 ;
        RECT 190.915 -33.485 191.245 -33.155 ;
        RECT 185.475 -33.485 185.805 -33.155 ;
        RECT 182.755 -33.485 183.085 -33.155 ;
        RECT 181.395 -33.485 181.725 -33.155 ;
        RECT 180.035 -33.485 180.365 -33.155 ;
        RECT 178.675 -33.485 179.005 -33.155 ;
        RECT 177.315 -33.485 177.645 -33.155 ;
        RECT 175.955 -33.485 176.285 -33.155 ;
        RECT 173.235 -33.485 173.565 -33.155 ;
        RECT 170.515 -33.485 170.845 -33.155 ;
        RECT 167.795 -33.485 168.125 -33.155 ;
        RECT 166.435 -33.485 166.765 -33.155 ;
        RECT 165.075 -33.485 165.405 -33.155 ;
        RECT 163.715 -33.485 164.045 -33.155 ;
        RECT 162.355 -33.485 162.685 -33.155 ;
        RECT 160.995 -33.485 161.325 -33.155 ;
        RECT 158.275 -33.485 158.605 -33.155 ;
        RECT 155.555 -33.485 155.885 -33.155 ;
        RECT 152.835 -33.485 153.165 -33.155 ;
        RECT 151.475 -33.485 151.805 -33.155 ;
        RECT 150.115 -33.485 150.445 -33.155 ;
        RECT 148.755 -33.485 149.085 -33.155 ;
        RECT 147.395 -33.485 147.725 -33.155 ;
        RECT 146.035 -33.485 146.365 -33.155 ;
        RECT 143.315 -33.485 143.645 -33.155 ;
        RECT 140.595 -33.485 140.925 -33.155 ;
        RECT 137.875 -33.485 138.205 -33.155 ;
        RECT 136.515 -33.485 136.845 -33.155 ;
        RECT 135.155 -33.485 135.485 -33.155 ;
        RECT 133.795 -33.485 134.125 -33.155 ;
        RECT 132.435 -33.485 132.765 -33.155 ;
        RECT 131.075 -33.485 131.405 -33.155 ;
        RECT 128.355 -33.485 128.685 -33.155 ;
        RECT 125.635 -33.485 125.965 -33.155 ;
        RECT 122.915 -33.485 123.245 -33.155 ;
        RECT 121.555 -33.485 121.885 -33.155 ;
        RECT 120.195 -33.485 120.525 -33.155 ;
        RECT 118.835 -33.485 119.165 -33.155 ;
        RECT 117.475 -33.485 117.805 -33.155 ;
        RECT 116.115 -33.485 116.445 -33.155 ;
        RECT 113.395 -33.485 113.725 -33.155 ;
        RECT 110.675 -33.485 111.005 -33.155 ;
        RECT 107.955 -33.485 108.285 -33.155 ;
        RECT 106.595 -33.485 106.925 -33.155 ;
        RECT 105.235 -33.485 105.565 -33.155 ;
        RECT 103.875 -33.485 104.205 -33.155 ;
        RECT 102.515 -33.485 102.845 -33.155 ;
        RECT 101.155 -33.485 101.485 -33.155 ;
        RECT 98.435 -33.485 98.765 -33.155 ;
        RECT 95.715 -33.485 96.045 -33.155 ;
        RECT 92.995 -33.485 93.325 -33.155 ;
        RECT 91.635 -33.485 91.965 -33.155 ;
        RECT 90.275 -33.485 90.605 -33.155 ;
        RECT 88.915 -33.485 89.245 -33.155 ;
        RECT 87.555 -33.485 87.885 -33.155 ;
        RECT 86.195 -33.485 86.525 -33.155 ;
        RECT 83.475 -33.485 83.805 -33.155 ;
        RECT 80.755 -33.485 81.085 -33.155 ;
        RECT 78.035 -33.485 78.365 -33.155 ;
        RECT 76.675 -33.485 77.005 -33.155 ;
        RECT 75.315 -33.485 75.645 -33.155 ;
        RECT 73.955 -33.485 74.285 -33.155 ;
        RECT 72.595 -33.485 72.925 -33.155 ;
        RECT 71.235 -33.485 71.565 -33.155 ;
        RECT 68.515 -33.485 68.845 -33.155 ;
        RECT 65.795 -33.485 66.125 -33.155 ;
        RECT 63.075 -33.485 63.405 -33.155 ;
        RECT 61.715 -33.485 62.045 -33.155 ;
        RECT 60.355 -33.485 60.685 -33.155 ;
        RECT 58.995 -33.485 59.325 -33.155 ;
        RECT 57.635 -33.485 57.965 -33.155 ;
        RECT 56.275 -33.485 56.605 -33.155 ;
        RECT 53.555 -33.485 53.885 -33.155 ;
        RECT 50.835 -33.485 51.165 -33.155 ;
        RECT 48.115 -33.485 48.445 -33.155 ;
        RECT 46.755 -33.485 47.085 -33.155 ;
        RECT 45.395 -33.485 45.725 -33.155 ;
        RECT 44.035 -33.485 44.365 -33.155 ;
        RECT 42.675 -33.485 43.005 -33.155 ;
        RECT 41.315 -33.485 41.645 -33.155 ;
        RECT 38.595 -33.485 38.925 -33.155 ;
        RECT 35.875 -33.485 36.205 -33.155 ;
        RECT 33.155 -33.485 33.485 -33.155 ;
        RECT 31.795 -33.485 32.125 -33.155 ;
        RECT 30.435 -33.485 30.765 -33.155 ;
        RECT 29.075 -33.485 29.405 -33.155 ;
        RECT 27.715 -33.485 28.045 -33.155 ;
        RECT 26.355 -33.485 26.685 -33.155 ;
        RECT 23.635 -33.485 23.965 -33.155 ;
        RECT 20.915 -33.485 21.245 -33.155 ;
        RECT 18.195 -33.485 18.525 -33.155 ;
        RECT 16.835 -33.485 17.165 -33.155 ;
        RECT 15.475 -33.485 15.805 -33.155 ;
        RECT 14.115 -33.485 14.445 -33.155 ;
        RECT 12.755 -33.485 13.085 -33.155 ;
        RECT 11.395 -33.485 11.725 -33.155 ;
        RECT 8.675 -33.485 9.005 -33.155 ;
        RECT 7.315 -33.485 7.645 -33.155 ;
        RECT 5.955 -33.485 6.285 -33.155 ;
        RECT 4.595 -33.485 4.925 -33.155 ;
        RECT 3.235 -33.485 3.565 -33.155 ;
        RECT 1.875 -33.485 2.205 -33.155 ;
        RECT 0.515 -33.485 0.845 -33.155 ;
        RECT -0.845 -33.485 -0.515 -33.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 949.12 -34.84 954.88 -34.52 ;
        RECT 953.875 -34.845 954.205 -34.515 ;
        RECT 952.515 -34.845 952.845 -34.515 ;
        RECT 951.155 -34.845 951.485 -34.515 ;
        RECT 949.795 -34.845 950.125 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -21.24 954.88 -20.92 ;
        RECT 953.875 -21.245 954.205 -20.915 ;
        RECT 952.515 -21.245 952.845 -20.915 ;
        RECT 951.155 -21.245 951.485 -20.915 ;
        RECT 949.795 -21.245 950.125 -20.915 ;
        RECT 947.075 -21.245 947.405 -20.915 ;
        RECT 945.715 -21.245 946.045 -20.915 ;
        RECT 942.995 -21.245 943.325 -20.915 ;
        RECT 940.275 -21.245 940.605 -20.915 ;
        RECT 938.915 -21.245 939.245 -20.915 ;
        RECT 937.555 -21.245 937.885 -20.915 ;
        RECT 936.195 -21.245 936.525 -20.915 ;
        RECT 934.835 -21.245 935.165 -20.915 ;
        RECT 932.115 -21.245 932.445 -20.915 ;
        RECT 930.755 -21.245 931.085 -20.915 ;
        RECT 928.035 -21.245 928.365 -20.915 ;
        RECT 925.315 -21.245 925.645 -20.915 ;
        RECT 923.955 -21.245 924.285 -20.915 ;
        RECT 922.595 -21.245 922.925 -20.915 ;
        RECT 921.235 -21.245 921.565 -20.915 ;
        RECT 919.875 -21.245 920.205 -20.915 ;
        RECT 917.155 -21.245 917.485 -20.915 ;
        RECT 913.075 -21.245 913.405 -20.915 ;
        RECT 910.355 -21.245 910.685 -20.915 ;
        RECT 908.995 -21.245 909.325 -20.915 ;
        RECT 907.635 -21.245 907.965 -20.915 ;
        RECT 906.275 -21.245 906.605 -20.915 ;
        RECT 904.915 -21.245 905.245 -20.915 ;
        RECT 902.195 -21.245 902.525 -20.915 ;
        RECT 898.115 -21.245 898.445 -20.915 ;
        RECT 895.395 -21.245 895.725 -20.915 ;
        RECT 894.035 -21.245 894.365 -20.915 ;
        RECT 892.675 -21.245 893.005 -20.915 ;
        RECT 891.315 -21.245 891.645 -20.915 ;
        RECT 889.955 -21.245 890.285 -20.915 ;
        RECT 887.235 -21.245 887.565 -20.915 ;
        RECT 883.155 -21.245 883.485 -20.915 ;
        RECT 880.435 -21.245 880.765 -20.915 ;
        RECT 879.075 -21.245 879.405 -20.915 ;
        RECT 877.715 -21.245 878.045 -20.915 ;
        RECT 876.355 -21.245 876.685 -20.915 ;
        RECT 874.995 -21.245 875.325 -20.915 ;
        RECT 872.275 -21.245 872.605 -20.915 ;
        RECT 868.195 -21.245 868.525 -20.915 ;
        RECT 865.475 -21.245 865.805 -20.915 ;
        RECT 864.115 -21.245 864.445 -20.915 ;
        RECT 862.755 -21.245 863.085 -20.915 ;
        RECT 861.395 -21.245 861.725 -20.915 ;
        RECT 860.035 -21.245 860.365 -20.915 ;
        RECT 857.315 -21.245 857.645 -20.915 ;
        RECT 853.235 -21.245 853.565 -20.915 ;
        RECT 850.515 -21.245 850.845 -20.915 ;
        RECT 849.155 -21.245 849.485 -20.915 ;
        RECT 847.795 -21.245 848.125 -20.915 ;
        RECT 846.435 -21.245 846.765 -20.915 ;
        RECT 843.715 -21.245 844.045 -20.915 ;
        RECT 842.355 -21.245 842.685 -20.915 ;
        RECT 838.275 -21.245 838.605 -20.915 ;
        RECT 835.555 -21.245 835.885 -20.915 ;
        RECT 834.195 -21.245 834.525 -20.915 ;
        RECT 832.835 -21.245 833.165 -20.915 ;
        RECT 831.475 -21.245 831.805 -20.915 ;
        RECT 828.755 -21.245 829.085 -20.915 ;
        RECT 827.395 -21.245 827.725 -20.915 ;
        RECT 823.315 -21.245 823.645 -20.915 ;
        RECT 820.595 -21.245 820.925 -20.915 ;
        RECT 819.235 -21.245 819.565 -20.915 ;
        RECT 817.875 -21.245 818.205 -20.915 ;
        RECT 816.515 -21.245 816.845 -20.915 ;
        RECT 813.795 -21.245 814.125 -20.915 ;
        RECT 812.435 -21.245 812.765 -20.915 ;
        RECT 806.995 -21.245 807.325 -20.915 ;
        RECT 805.635 -21.245 805.965 -20.915 ;
        RECT 804.275 -21.245 804.605 -20.915 ;
        RECT 802.915 -21.245 803.245 -20.915 ;
        RECT 801.555 -21.245 801.885 -20.915 ;
        RECT 798.835 -21.245 799.165 -20.915 ;
        RECT 797.475 -21.245 797.805 -20.915 ;
        RECT 792.035 -21.245 792.365 -20.915 ;
        RECT 790.675 -21.245 791.005 -20.915 ;
        RECT 789.315 -21.245 789.645 -20.915 ;
        RECT 787.955 -21.245 788.285 -20.915 ;
        RECT 786.595 -21.245 786.925 -20.915 ;
        RECT 783.875 -21.245 784.205 -20.915 ;
        RECT 782.515 -21.245 782.845 -20.915 ;
        RECT 777.075 -21.245 777.405 -20.915 ;
        RECT 775.715 -21.245 776.045 -20.915 ;
        RECT 774.355 -21.245 774.685 -20.915 ;
        RECT 772.995 -21.245 773.325 -20.915 ;
        RECT 771.635 -21.245 771.965 -20.915 ;
        RECT 768.915 -21.245 769.245 -20.915 ;
        RECT 767.555 -21.245 767.885 -20.915 ;
        RECT 762.115 -21.245 762.445 -20.915 ;
        RECT 760.755 -21.245 761.085 -20.915 ;
        RECT 759.395 -21.245 759.725 -20.915 ;
        RECT 758.035 -21.245 758.365 -20.915 ;
        RECT 756.675 -21.245 757.005 -20.915 ;
        RECT 753.955 -21.245 754.285 -20.915 ;
        RECT 752.595 -21.245 752.925 -20.915 ;
        RECT 747.155 -21.245 747.485 -20.915 ;
        RECT 745.795 -21.245 746.125 -20.915 ;
        RECT 744.435 -21.245 744.765 -20.915 ;
        RECT 743.075 -21.245 743.405 -20.915 ;
        RECT 741.715 -21.245 742.045 -20.915 ;
        RECT 738.995 -21.245 739.325 -20.915 ;
        RECT 737.635 -21.245 737.965 -20.915 ;
        RECT 732.195 -21.245 732.525 -20.915 ;
        RECT 730.835 -21.245 731.165 -20.915 ;
        RECT 729.475 -21.245 729.805 -20.915 ;
        RECT 728.115 -21.245 728.445 -20.915 ;
        RECT 726.755 -21.245 727.085 -20.915 ;
        RECT 724.035 -21.245 724.365 -20.915 ;
        RECT 722.675 -21.245 723.005 -20.915 ;
        RECT 717.235 -21.245 717.565 -20.915 ;
        RECT 715.875 -21.245 716.205 -20.915 ;
        RECT 714.515 -21.245 714.845 -20.915 ;
        RECT 713.155 -21.245 713.485 -20.915 ;
        RECT 711.795 -21.245 712.125 -20.915 ;
        RECT 709.075 -21.245 709.405 -20.915 ;
        RECT 707.715 -21.245 708.045 -20.915 ;
        RECT 702.275 -21.245 702.605 -20.915 ;
        RECT 700.915 -21.245 701.245 -20.915 ;
        RECT 699.555 -21.245 699.885 -20.915 ;
        RECT 698.195 -21.245 698.525 -20.915 ;
        RECT 696.835 -21.245 697.165 -20.915 ;
        RECT 694.115 -21.245 694.445 -20.915 ;
        RECT 692.755 -21.245 693.085 -20.915 ;
        RECT 687.315 -21.245 687.645 -20.915 ;
        RECT 685.955 -21.245 686.285 -20.915 ;
        RECT 684.595 -21.245 684.925 -20.915 ;
        RECT 683.235 -21.245 683.565 -20.915 ;
        RECT 681.875 -21.245 682.205 -20.915 ;
        RECT 679.155 -21.245 679.485 -20.915 ;
        RECT 677.795 -21.245 678.125 -20.915 ;
        RECT 672.355 -21.245 672.685 -20.915 ;
        RECT 670.995 -21.245 671.325 -20.915 ;
        RECT 669.635 -21.245 669.965 -20.915 ;
        RECT 668.275 -21.245 668.605 -20.915 ;
        RECT 666.915 -21.245 667.245 -20.915 ;
        RECT 664.195 -21.245 664.525 -20.915 ;
        RECT 662.835 -21.245 663.165 -20.915 ;
        RECT 657.395 -21.245 657.725 -20.915 ;
        RECT 656.035 -21.245 656.365 -20.915 ;
        RECT 654.675 -21.245 655.005 -20.915 ;
        RECT 653.315 -21.245 653.645 -20.915 ;
        RECT 651.955 -21.245 652.285 -20.915 ;
        RECT 649.235 -21.245 649.565 -20.915 ;
        RECT 647.875 -21.245 648.205 -20.915 ;
        RECT 642.435 -21.245 642.765 -20.915 ;
        RECT 641.075 -21.245 641.405 -20.915 ;
        RECT 639.715 -21.245 640.045 -20.915 ;
        RECT 638.355 -21.245 638.685 -20.915 ;
        RECT 636.995 -21.245 637.325 -20.915 ;
        RECT 634.275 -21.245 634.605 -20.915 ;
        RECT 632.915 -21.245 633.245 -20.915 ;
        RECT 627.475 -21.245 627.805 -20.915 ;
        RECT 626.115 -21.245 626.445 -20.915 ;
        RECT 624.755 -21.245 625.085 -20.915 ;
        RECT 623.395 -21.245 623.725 -20.915 ;
        RECT 622.035 -21.245 622.365 -20.915 ;
        RECT 619.315 -21.245 619.645 -20.915 ;
        RECT 617.955 -21.245 618.285 -20.915 ;
        RECT 612.515 -21.245 612.845 -20.915 ;
        RECT 611.155 -21.245 611.485 -20.915 ;
        RECT 609.795 -21.245 610.125 -20.915 ;
        RECT 608.435 -21.245 608.765 -20.915 ;
        RECT 607.075 -21.245 607.405 -20.915 ;
        RECT 604.355 -21.245 604.685 -20.915 ;
        RECT 602.995 -21.245 603.325 -20.915 ;
        RECT 600.275 -21.245 600.605 -20.915 ;
        RECT 597.555 -21.245 597.885 -20.915 ;
        RECT 596.195 -21.245 596.525 -20.915 ;
        RECT 594.835 -21.245 595.165 -20.915 ;
        RECT 593.475 -21.245 593.805 -20.915 ;
        RECT 592.115 -21.245 592.445 -20.915 ;
        RECT 589.395 -21.245 589.725 -20.915 ;
        RECT 588.035 -21.245 588.365 -20.915 ;
        RECT 585.315 -21.245 585.645 -20.915 ;
        RECT 582.595 -21.245 582.925 -20.915 ;
        RECT 581.235 -21.245 581.565 -20.915 ;
        RECT 579.875 -21.245 580.205 -20.915 ;
        RECT 578.515 -21.245 578.845 -20.915 ;
        RECT 577.155 -21.245 577.485 -20.915 ;
        RECT 574.435 -21.245 574.765 -20.915 ;
        RECT 570.355 -21.245 570.685 -20.915 ;
        RECT 567.635 -21.245 567.965 -20.915 ;
        RECT 566.275 -21.245 566.605 -20.915 ;
        RECT 564.915 -21.245 565.245 -20.915 ;
        RECT 563.555 -21.245 563.885 -20.915 ;
        RECT 562.195 -21.245 562.525 -20.915 ;
        RECT 559.475 -21.245 559.805 -20.915 ;
        RECT 555.395 -21.245 555.725 -20.915 ;
        RECT 552.675 -21.245 553.005 -20.915 ;
        RECT 551.315 -21.245 551.645 -20.915 ;
        RECT 549.955 -21.245 550.285 -20.915 ;
        RECT 548.595 -21.245 548.925 -20.915 ;
        RECT 547.235 -21.245 547.565 -20.915 ;
        RECT 544.515 -21.245 544.845 -20.915 ;
        RECT 540.435 -21.245 540.765 -20.915 ;
        RECT 537.715 -21.245 538.045 -20.915 ;
        RECT 536.355 -21.245 536.685 -20.915 ;
        RECT 534.995 -21.245 535.325 -20.915 ;
        RECT 533.635 -21.245 533.965 -20.915 ;
        RECT 532.275 -21.245 532.605 -20.915 ;
        RECT 529.555 -21.245 529.885 -20.915 ;
        RECT 525.475 -21.245 525.805 -20.915 ;
        RECT 522.755 -21.245 523.085 -20.915 ;
        RECT 521.395 -21.245 521.725 -20.915 ;
        RECT 520.035 -21.245 520.365 -20.915 ;
        RECT 518.675 -21.245 519.005 -20.915 ;
        RECT 517.315 -21.245 517.645 -20.915 ;
        RECT 515.955 -21.245 516.285 -20.915 ;
        RECT 514.595 -21.245 514.925 -20.915 ;
        RECT 510.515 -21.245 510.845 -20.915 ;
        RECT 507.795 -21.245 508.125 -20.915 ;
        RECT 506.435 -21.245 506.765 -20.915 ;
        RECT 505.075 -21.245 505.405 -20.915 ;
        RECT 503.715 -21.245 504.045 -20.915 ;
        RECT 500.995 -21.245 501.325 -20.915 ;
        RECT 499.635 -21.245 499.965 -20.915 ;
        RECT 495.555 -21.245 495.885 -20.915 ;
        RECT 492.835 -21.245 493.165 -20.915 ;
        RECT 491.475 -21.245 491.805 -20.915 ;
        RECT 490.115 -21.245 490.445 -20.915 ;
        RECT 488.755 -21.245 489.085 -20.915 ;
        RECT 486.035 -21.245 486.365 -20.915 ;
        RECT 484.675 -21.245 485.005 -20.915 ;
        RECT 480.595 -21.245 480.925 -20.915 ;
        RECT 477.875 -21.245 478.205 -20.915 ;
        RECT 476.515 -21.245 476.845 -20.915 ;
        RECT 475.155 -21.245 475.485 -20.915 ;
        RECT 473.795 -21.245 474.125 -20.915 ;
        RECT 471.075 -21.245 471.405 -20.915 ;
        RECT 469.715 -21.245 470.045 -20.915 ;
        RECT 464.275 -21.245 464.605 -20.915 ;
        RECT 462.915 -21.245 463.245 -20.915 ;
        RECT 461.555 -21.245 461.885 -20.915 ;
        RECT 460.195 -21.245 460.525 -20.915 ;
        RECT 458.835 -21.245 459.165 -20.915 ;
        RECT 456.115 -21.245 456.445 -20.915 ;
        RECT 454.755 -21.245 455.085 -20.915 ;
        RECT 449.315 -21.245 449.645 -20.915 ;
        RECT 447.955 -21.245 448.285 -20.915 ;
        RECT 446.595 -21.245 446.925 -20.915 ;
        RECT 445.235 -21.245 445.565 -20.915 ;
        RECT 443.875 -21.245 444.205 -20.915 ;
        RECT 441.155 -21.245 441.485 -20.915 ;
        RECT 439.795 -21.245 440.125 -20.915 ;
        RECT 434.355 -21.245 434.685 -20.915 ;
        RECT 432.995 -21.245 433.325 -20.915 ;
        RECT 431.635 -21.245 431.965 -20.915 ;
        RECT 430.275 -21.245 430.605 -20.915 ;
        RECT 428.915 -21.245 429.245 -20.915 ;
        RECT 426.195 -21.245 426.525 -20.915 ;
        RECT 424.835 -21.245 425.165 -20.915 ;
        RECT 419.395 -21.245 419.725 -20.915 ;
        RECT 418.035 -21.245 418.365 -20.915 ;
        RECT 416.675 -21.245 417.005 -20.915 ;
        RECT 415.315 -21.245 415.645 -20.915 ;
        RECT 413.955 -21.245 414.285 -20.915 ;
        RECT 411.235 -21.245 411.565 -20.915 ;
        RECT 409.875 -21.245 410.205 -20.915 ;
        RECT 404.435 -21.245 404.765 -20.915 ;
        RECT 403.075 -21.245 403.405 -20.915 ;
        RECT 401.715 -21.245 402.045 -20.915 ;
        RECT 400.355 -21.245 400.685 -20.915 ;
        RECT 398.995 -21.245 399.325 -20.915 ;
        RECT 396.275 -21.245 396.605 -20.915 ;
        RECT 394.915 -21.245 395.245 -20.915 ;
        RECT 389.475 -21.245 389.805 -20.915 ;
        RECT 388.115 -21.245 388.445 -20.915 ;
        RECT 386.755 -21.245 387.085 -20.915 ;
        RECT 385.395 -21.245 385.725 -20.915 ;
        RECT 384.035 -21.245 384.365 -20.915 ;
        RECT 381.315 -21.245 381.645 -20.915 ;
        RECT 379.955 -21.245 380.285 -20.915 ;
        RECT 374.515 -21.245 374.845 -20.915 ;
        RECT 373.155 -21.245 373.485 -20.915 ;
        RECT 371.795 -21.245 372.125 -20.915 ;
        RECT 370.435 -21.245 370.765 -20.915 ;
        RECT 369.075 -21.245 369.405 -20.915 ;
        RECT 366.355 -21.245 366.685 -20.915 ;
        RECT 364.995 -21.245 365.325 -20.915 ;
        RECT 359.555 -21.245 359.885 -20.915 ;
        RECT 358.195 -21.245 358.525 -20.915 ;
        RECT 356.835 -21.245 357.165 -20.915 ;
        RECT 355.475 -21.245 355.805 -20.915 ;
        RECT 354.115 -21.245 354.445 -20.915 ;
        RECT 351.395 -21.245 351.725 -20.915 ;
        RECT 350.035 -21.245 350.365 -20.915 ;
        RECT 344.595 -21.245 344.925 -20.915 ;
        RECT 343.235 -21.245 343.565 -20.915 ;
        RECT 341.875 -21.245 342.205 -20.915 ;
        RECT 340.515 -21.245 340.845 -20.915 ;
        RECT 339.155 -21.245 339.485 -20.915 ;
        RECT 336.435 -21.245 336.765 -20.915 ;
        RECT 335.075 -21.245 335.405 -20.915 ;
        RECT 329.635 -21.245 329.965 -20.915 ;
        RECT 328.275 -21.245 328.605 -20.915 ;
        RECT 326.915 -21.245 327.245 -20.915 ;
        RECT 325.555 -21.245 325.885 -20.915 ;
        RECT 324.195 -21.245 324.525 -20.915 ;
        RECT 321.475 -21.245 321.805 -20.915 ;
        RECT 320.115 -21.245 320.445 -20.915 ;
        RECT 314.675 -21.245 315.005 -20.915 ;
        RECT 313.315 -21.245 313.645 -20.915 ;
        RECT 311.955 -21.245 312.285 -20.915 ;
        RECT 310.595 -21.245 310.925 -20.915 ;
        RECT 309.235 -21.245 309.565 -20.915 ;
        RECT 306.515 -21.245 306.845 -20.915 ;
        RECT 305.155 -21.245 305.485 -20.915 ;
        RECT 299.715 -21.245 300.045 -20.915 ;
        RECT 298.355 -21.245 298.685 -20.915 ;
        RECT 296.995 -21.245 297.325 -20.915 ;
        RECT 295.635 -21.245 295.965 -20.915 ;
        RECT 294.275 -21.245 294.605 -20.915 ;
        RECT 291.555 -21.245 291.885 -20.915 ;
        RECT 290.195 -21.245 290.525 -20.915 ;
        RECT 284.755 -21.245 285.085 -20.915 ;
        RECT 283.395 -21.245 283.725 -20.915 ;
        RECT 282.035 -21.245 282.365 -20.915 ;
        RECT 280.675 -21.245 281.005 -20.915 ;
        RECT 279.315 -21.245 279.645 -20.915 ;
        RECT 276.595 -21.245 276.925 -20.915 ;
        RECT 275.235 -21.245 275.565 -20.915 ;
        RECT 272.515 -21.245 272.845 -20.915 ;
        RECT 269.795 -21.245 270.125 -20.915 ;
        RECT 268.435 -21.245 268.765 -20.915 ;
        RECT 267.075 -21.245 267.405 -20.915 ;
        RECT 265.715 -21.245 266.045 -20.915 ;
        RECT 264.355 -21.245 264.685 -20.915 ;
        RECT 261.635 -21.245 261.965 -20.915 ;
        RECT 260.275 -21.245 260.605 -20.915 ;
        RECT 257.555 -21.245 257.885 -20.915 ;
        RECT 254.835 -21.245 255.165 -20.915 ;
        RECT 253.475 -21.245 253.805 -20.915 ;
        RECT 252.115 -21.245 252.445 -20.915 ;
        RECT 250.755 -21.245 251.085 -20.915 ;
        RECT 249.395 -21.245 249.725 -20.915 ;
        RECT 246.675 -21.245 247.005 -20.915 ;
        RECT 242.595 -21.245 242.925 -20.915 ;
        RECT 239.875 -21.245 240.205 -20.915 ;
        RECT 238.515 -21.245 238.845 -20.915 ;
        RECT 237.155 -21.245 237.485 -20.915 ;
        RECT 235.795 -21.245 236.125 -20.915 ;
        RECT 234.435 -21.245 234.765 -20.915 ;
        RECT 231.715 -21.245 232.045 -20.915 ;
        RECT 227.635 -21.245 227.965 -20.915 ;
        RECT 224.915 -21.245 225.245 -20.915 ;
        RECT 223.555 -21.245 223.885 -20.915 ;
        RECT 222.195 -21.245 222.525 -20.915 ;
        RECT 220.835 -21.245 221.165 -20.915 ;
        RECT 219.475 -21.245 219.805 -20.915 ;
        RECT 216.755 -21.245 217.085 -20.915 ;
        RECT 212.675 -21.245 213.005 -20.915 ;
        RECT 209.955 -21.245 210.285 -20.915 ;
        RECT 208.595 -21.245 208.925 -20.915 ;
        RECT 207.235 -21.245 207.565 -20.915 ;
        RECT 205.875 -21.245 206.205 -20.915 ;
        RECT 204.515 -21.245 204.845 -20.915 ;
        RECT 201.795 -21.245 202.125 -20.915 ;
        RECT 197.715 -21.245 198.045 -20.915 ;
        RECT 194.995 -21.245 195.325 -20.915 ;
        RECT 193.635 -21.245 193.965 -20.915 ;
        RECT 192.275 -21.245 192.605 -20.915 ;
        RECT 190.915 -21.245 191.245 -20.915 ;
        RECT 189.555 -21.245 189.885 -20.915 ;
        RECT 186.835 -21.245 187.165 -20.915 ;
        RECT 182.755 -21.245 183.085 -20.915 ;
        RECT 180.035 -21.245 180.365 -20.915 ;
        RECT 178.675 -21.245 179.005 -20.915 ;
        RECT 177.315 -21.245 177.645 -20.915 ;
        RECT 175.955 -21.245 176.285 -20.915 ;
        RECT 173.235 -21.245 173.565 -20.915 ;
        RECT 171.875 -21.245 172.205 -20.915 ;
        RECT 167.795 -21.245 168.125 -20.915 ;
        RECT 165.075 -21.245 165.405 -20.915 ;
        RECT 163.715 -21.245 164.045 -20.915 ;
        RECT 162.355 -21.245 162.685 -20.915 ;
        RECT 160.995 -21.245 161.325 -20.915 ;
        RECT 158.275 -21.245 158.605 -20.915 ;
        RECT 156.915 -21.245 157.245 -20.915 ;
        RECT 152.835 -21.245 153.165 -20.915 ;
        RECT 150.115 -21.245 150.445 -20.915 ;
        RECT 148.755 -21.245 149.085 -20.915 ;
        RECT 147.395 -21.245 147.725 -20.915 ;
        RECT 146.035 -21.245 146.365 -20.915 ;
        RECT 143.315 -21.245 143.645 -20.915 ;
        RECT 141.955 -21.245 142.285 -20.915 ;
        RECT 136.515 -21.245 136.845 -20.915 ;
        RECT 135.155 -21.245 135.485 -20.915 ;
        RECT 133.795 -21.245 134.125 -20.915 ;
        RECT 132.435 -21.245 132.765 -20.915 ;
        RECT 131.075 -21.245 131.405 -20.915 ;
        RECT 128.355 -21.245 128.685 -20.915 ;
        RECT 126.995 -21.245 127.325 -20.915 ;
        RECT 121.555 -21.245 121.885 -20.915 ;
        RECT 120.195 -21.245 120.525 -20.915 ;
        RECT 118.835 -21.245 119.165 -20.915 ;
        RECT 117.475 -21.245 117.805 -20.915 ;
        RECT 116.115 -21.245 116.445 -20.915 ;
        RECT 113.395 -21.245 113.725 -20.915 ;
        RECT 112.035 -21.245 112.365 -20.915 ;
        RECT 106.595 -21.245 106.925 -20.915 ;
        RECT 105.235 -21.245 105.565 -20.915 ;
        RECT 103.875 -21.245 104.205 -20.915 ;
        RECT 102.515 -21.245 102.845 -20.915 ;
        RECT 101.155 -21.245 101.485 -20.915 ;
        RECT 98.435 -21.245 98.765 -20.915 ;
        RECT 97.075 -21.245 97.405 -20.915 ;
        RECT 91.635 -21.245 91.965 -20.915 ;
        RECT 90.275 -21.245 90.605 -20.915 ;
        RECT 88.915 -21.245 89.245 -20.915 ;
        RECT 87.555 -21.245 87.885 -20.915 ;
        RECT 86.195 -21.245 86.525 -20.915 ;
        RECT 83.475 -21.245 83.805 -20.915 ;
        RECT 82.115 -21.245 82.445 -20.915 ;
        RECT 76.675 -21.245 77.005 -20.915 ;
        RECT 75.315 -21.245 75.645 -20.915 ;
        RECT 73.955 -21.245 74.285 -20.915 ;
        RECT 72.595 -21.245 72.925 -20.915 ;
        RECT 71.235 -21.245 71.565 -20.915 ;
        RECT 68.515 -21.245 68.845 -20.915 ;
        RECT 67.155 -21.245 67.485 -20.915 ;
        RECT 61.715 -21.245 62.045 -20.915 ;
        RECT 60.355 -21.245 60.685 -20.915 ;
        RECT 58.995 -21.245 59.325 -20.915 ;
        RECT 57.635 -21.245 57.965 -20.915 ;
        RECT 56.275 -21.245 56.605 -20.915 ;
        RECT 53.555 -21.245 53.885 -20.915 ;
        RECT 52.195 -21.245 52.525 -20.915 ;
        RECT 46.755 -21.245 47.085 -20.915 ;
        RECT 45.395 -21.245 45.725 -20.915 ;
        RECT 44.035 -21.245 44.365 -20.915 ;
        RECT 42.675 -21.245 43.005 -20.915 ;
        RECT 41.315 -21.245 41.645 -20.915 ;
        RECT 38.595 -21.245 38.925 -20.915 ;
        RECT 37.235 -21.245 37.565 -20.915 ;
        RECT 31.795 -21.245 32.125 -20.915 ;
        RECT 30.435 -21.245 30.765 -20.915 ;
        RECT 29.075 -21.245 29.405 -20.915 ;
        RECT 27.715 -21.245 28.045 -20.915 ;
        RECT 26.355 -21.245 26.685 -20.915 ;
        RECT 23.635 -21.245 23.965 -20.915 ;
        RECT 22.275 -21.245 22.605 -20.915 ;
        RECT 16.835 -21.245 17.165 -20.915 ;
        RECT 15.475 -21.245 15.805 -20.915 ;
        RECT 14.115 -21.245 14.445 -20.915 ;
        RECT 12.755 -21.245 13.085 -20.915 ;
        RECT 11.395 -21.245 11.725 -20.915 ;
        RECT 8.675 -21.245 9.005 -20.915 ;
        RECT 7.315 -21.245 7.645 -20.915 ;
        RECT 3.235 -21.245 3.565 -20.915 ;
        RECT 1.875 -21.245 2.205 -20.915 ;
        RECT 0.515 -21.245 0.845 -20.915 ;
        RECT -0.845 -21.245 -0.515 -20.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 943.68 -23.96 954.88 -23.64 ;
        RECT 953.875 -23.965 954.205 -23.635 ;
        RECT 952.515 -23.965 952.845 -23.635 ;
        RECT 951.155 -23.965 951.485 -23.635 ;
        RECT 949.795 -23.965 950.125 -23.635 ;
        RECT 947.075 -23.965 947.405 -23.635 ;
        RECT 945.715 -23.965 946.045 -23.635 ;
        RECT 944.355 -23.965 944.685 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 934.84 -26.68 954.88 -26.36 ;
        RECT 953.875 -26.685 954.205 -26.355 ;
        RECT 952.515 -26.685 952.845 -26.355 ;
        RECT 951.155 -26.685 951.485 -26.355 ;
        RECT 949.795 -26.685 950.125 -26.355 ;
        RECT 947.075 -26.685 947.405 -26.355 ;
        RECT 945.715 -26.685 946.045 -26.355 ;
        RECT 944.355 -26.685 944.685 -26.355 ;
        RECT 942.995 -26.685 943.325 -26.355 ;
        RECT 941.635 -26.685 941.965 -26.355 ;
        RECT 940.275 -26.685 940.605 -26.355 ;
        RECT 938.915 -26.685 939.245 -26.355 ;
        RECT 937.555 -26.685 937.885 -26.355 ;
        RECT 936.195 -26.685 936.525 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 930.76 -28.04 954.88 -27.72 ;
        RECT 953.875 -28.045 954.205 -27.715 ;
        RECT 952.515 -28.045 952.845 -27.715 ;
        RECT 951.155 -28.045 951.485 -27.715 ;
        RECT 949.795 -28.045 950.125 -27.715 ;
        RECT 947.075 -28.045 947.405 -27.715 ;
        RECT 945.715 -28.045 946.045 -27.715 ;
        RECT 944.355 -28.045 944.685 -27.715 ;
        RECT 942.995 -28.045 943.325 -27.715 ;
        RECT 941.635 -28.045 941.965 -27.715 ;
        RECT 940.275 -28.045 940.605 -27.715 ;
        RECT 938.915 -28.045 939.245 -27.715 ;
        RECT 937.555 -28.045 937.885 -27.715 ;
        RECT 936.195 -28.045 936.525 -27.715 ;
        RECT 932.115 -28.045 932.445 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 934.84 -29.4 954.88 -29.08 ;
        RECT 953.875 -29.405 954.205 -29.075 ;
        RECT 952.515 -29.405 952.845 -29.075 ;
        RECT 951.155 -29.405 951.485 -29.075 ;
        RECT 949.795 -29.405 950.125 -29.075 ;
        RECT 947.075 -29.405 947.405 -29.075 ;
        RECT 945.715 -29.405 946.045 -29.075 ;
        RECT 944.355 -29.405 944.685 -29.075 ;
        RECT 942.995 -29.405 943.325 -29.075 ;
        RECT 941.635 -29.405 941.965 -29.075 ;
        RECT 940.275 -29.405 940.605 -29.075 ;
        RECT 938.915 -29.405 939.245 -29.075 ;
        RECT 937.555 -29.405 937.885 -29.075 ;
        RECT 936.195 -29.405 936.525 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 938.915 -30.765 939.245 -30.435 ;
        RECT 937.555 -30.765 937.885 -30.435 ;
        RECT 936.195 -30.765 936.525 -30.435 ;
        RECT 932.115 -30.765 932.445 -30.435 ;
        RECT 928.035 -30.765 928.365 -30.435 ;
        RECT 925.315 -30.765 925.645 -30.435 ;
        RECT 923.955 -30.765 924.285 -30.435 ;
        RECT 922.595 -30.765 922.925 -30.435 ;
        RECT 921.235 -30.765 921.565 -30.435 ;
        RECT 917.155 -30.765 917.485 -30.435 ;
        RECT 913.075 -30.765 913.405 -30.435 ;
        RECT 910.355 -30.765 910.685 -30.435 ;
        RECT 908.995 -30.765 909.325 -30.435 ;
        RECT 907.635 -30.765 907.965 -30.435 ;
        RECT 906.275 -30.765 906.605 -30.435 ;
        RECT 902.195 -30.765 902.525 -30.435 ;
        RECT 900.835 -30.765 901.165 -30.435 ;
        RECT 898.115 -30.765 898.445 -30.435 ;
        RECT 895.395 -30.765 895.725 -30.435 ;
        RECT 894.035 -30.765 894.365 -30.435 ;
        RECT 892.675 -30.765 893.005 -30.435 ;
        RECT 891.315 -30.765 891.645 -30.435 ;
        RECT 885.875 -30.765 886.205 -30.435 ;
        RECT 883.155 -30.765 883.485 -30.435 ;
        RECT 880.435 -30.765 880.765 -30.435 ;
        RECT 879.075 -30.765 879.405 -30.435 ;
        RECT 877.715 -30.765 878.045 -30.435 ;
        RECT 876.355 -30.765 876.685 -30.435 ;
        RECT 870.915 -30.765 871.245 -30.435 ;
        RECT 868.195 -30.765 868.525 -30.435 ;
        RECT 865.475 -30.765 865.805 -30.435 ;
        RECT 864.115 -30.765 864.445 -30.435 ;
        RECT 862.755 -30.765 863.085 -30.435 ;
        RECT 861.395 -30.765 861.725 -30.435 ;
        RECT 855.955 -30.765 856.285 -30.435 ;
        RECT 853.235 -30.765 853.565 -30.435 ;
        RECT 850.515 -30.765 850.845 -30.435 ;
        RECT 849.155 -30.765 849.485 -30.435 ;
        RECT 847.795 -30.765 848.125 -30.435 ;
        RECT 846.435 -30.765 846.765 -30.435 ;
        RECT 840.995 -30.765 841.325 -30.435 ;
        RECT 838.275 -30.765 838.605 -30.435 ;
        RECT 835.555 -30.765 835.885 -30.435 ;
        RECT 834.195 -30.765 834.525 -30.435 ;
        RECT 832.835 -30.765 833.165 -30.435 ;
        RECT 831.475 -30.765 831.805 -30.435 ;
        RECT 826.035 -30.765 826.365 -30.435 ;
        RECT 823.315 -30.765 823.645 -30.435 ;
        RECT 820.595 -30.765 820.925 -30.435 ;
        RECT 819.235 -30.765 819.565 -30.435 ;
        RECT 817.875 -30.765 818.205 -30.435 ;
        RECT 816.515 -30.765 816.845 -30.435 ;
        RECT 811.075 -30.765 811.405 -30.435 ;
        RECT 808.355 -30.765 808.685 -30.435 ;
        RECT 805.635 -30.765 805.965 -30.435 ;
        RECT 804.275 -30.765 804.605 -30.435 ;
        RECT 802.915 -30.765 803.245 -30.435 ;
        RECT 801.555 -30.765 801.885 -30.435 ;
        RECT 796.115 -30.765 796.445 -30.435 ;
        RECT 793.395 -30.765 793.725 -30.435 ;
        RECT 790.675 -30.765 791.005 -30.435 ;
        RECT 789.315 -30.765 789.645 -30.435 ;
        RECT 787.955 -30.765 788.285 -30.435 ;
        RECT 786.595 -30.765 786.925 -30.435 ;
        RECT 781.155 -30.765 781.485 -30.435 ;
        RECT 778.435 -30.765 778.765 -30.435 ;
        RECT 775.715 -30.765 776.045 -30.435 ;
        RECT 774.355 -30.765 774.685 -30.435 ;
        RECT 772.995 -30.765 773.325 -30.435 ;
        RECT 771.635 -30.765 771.965 -30.435 ;
        RECT 766.195 -30.765 766.525 -30.435 ;
        RECT 763.475 -30.765 763.805 -30.435 ;
        RECT 760.755 -30.765 761.085 -30.435 ;
        RECT 759.395 -30.765 759.725 -30.435 ;
        RECT 758.035 -30.765 758.365 -30.435 ;
        RECT 756.675 -30.765 757.005 -30.435 ;
        RECT 751.235 -30.765 751.565 -30.435 ;
        RECT 748.515 -30.765 748.845 -30.435 ;
        RECT 745.795 -30.765 746.125 -30.435 ;
        RECT 744.435 -30.765 744.765 -30.435 ;
        RECT 743.075 -30.765 743.405 -30.435 ;
        RECT 741.715 -30.765 742.045 -30.435 ;
        RECT 736.275 -30.765 736.605 -30.435 ;
        RECT 733.555 -30.765 733.885 -30.435 ;
        RECT 730.835 -30.765 731.165 -30.435 ;
        RECT 729.475 -30.765 729.805 -30.435 ;
        RECT 728.115 -30.765 728.445 -30.435 ;
        RECT 726.755 -30.765 727.085 -30.435 ;
        RECT 721.315 -30.765 721.645 -30.435 ;
        RECT 718.595 -30.765 718.925 -30.435 ;
        RECT 715.875 -30.765 716.205 -30.435 ;
        RECT 714.515 -30.765 714.845 -30.435 ;
        RECT 713.155 -30.765 713.485 -30.435 ;
        RECT 711.795 -30.765 712.125 -30.435 ;
        RECT 706.355 -30.765 706.685 -30.435 ;
        RECT 703.635 -30.765 703.965 -30.435 ;
        RECT 700.915 -30.765 701.245 -30.435 ;
        RECT 699.555 -30.765 699.885 -30.435 ;
        RECT 698.195 -30.765 698.525 -30.435 ;
        RECT 696.835 -30.765 697.165 -30.435 ;
        RECT 691.395 -30.765 691.725 -30.435 ;
        RECT 688.675 -30.765 689.005 -30.435 ;
        RECT 685.955 -30.765 686.285 -30.435 ;
        RECT 684.595 -30.765 684.925 -30.435 ;
        RECT 683.235 -30.765 683.565 -30.435 ;
        RECT 681.875 -30.765 682.205 -30.435 ;
        RECT 679.155 -30.765 679.485 -30.435 ;
        RECT 676.435 -30.765 676.765 -30.435 ;
        RECT 673.715 -30.765 674.045 -30.435 ;
        RECT 670.995 -30.765 671.325 -30.435 ;
        RECT 669.635 -30.765 669.965 -30.435 ;
        RECT 668.275 -30.765 668.605 -30.435 ;
        RECT 664.195 -30.765 664.525 -30.435 ;
        RECT 661.475 -30.765 661.805 -30.435 ;
        RECT 658.755 -30.765 659.085 -30.435 ;
        RECT 656.035 -30.765 656.365 -30.435 ;
        RECT 654.675 -30.765 655.005 -30.435 ;
        RECT 653.315 -30.765 653.645 -30.435 ;
        RECT 649.235 -30.765 649.565 -30.435 ;
        RECT 646.515 -30.765 646.845 -30.435 ;
        RECT 643.795 -30.765 644.125 -30.435 ;
        RECT 641.075 -30.765 641.405 -30.435 ;
        RECT 639.715 -30.765 640.045 -30.435 ;
        RECT 638.355 -30.765 638.685 -30.435 ;
        RECT 634.275 -30.765 634.605 -30.435 ;
        RECT 631.555 -30.765 631.885 -30.435 ;
        RECT 627.475 -30.765 627.805 -30.435 ;
        RECT 626.115 -30.765 626.445 -30.435 ;
        RECT 624.755 -30.765 625.085 -30.435 ;
        RECT 623.395 -30.765 623.725 -30.435 ;
        RECT 619.315 -30.765 619.645 -30.435 ;
        RECT 616.595 -30.765 616.925 -30.435 ;
        RECT 612.515 -30.765 612.845 -30.435 ;
        RECT 611.155 -30.765 611.485 -30.435 ;
        RECT 609.795 -30.765 610.125 -30.435 ;
        RECT 608.435 -30.765 608.765 -30.435 ;
        RECT 604.355 -30.765 604.685 -30.435 ;
        RECT 600.275 -30.765 600.605 -30.435 ;
        RECT 597.555 -30.765 597.885 -30.435 ;
        RECT 596.195 -30.765 596.525 -30.435 ;
        RECT 594.835 -30.765 595.165 -30.435 ;
        RECT 593.475 -30.765 593.805 -30.435 ;
        RECT 589.395 -30.765 589.725 -30.435 ;
        RECT 585.315 -30.765 585.645 -30.435 ;
        RECT 582.595 -30.765 582.925 -30.435 ;
        RECT 581.235 -30.765 581.565 -30.435 ;
        RECT 579.875 -30.765 580.205 -30.435 ;
        RECT 578.515 -30.765 578.845 -30.435 ;
        RECT 574.435 -30.765 574.765 -30.435 ;
        RECT 570.355 -30.765 570.685 -30.435 ;
        RECT 567.635 -30.765 567.965 -30.435 ;
        RECT 566.275 -30.765 566.605 -30.435 ;
        RECT 564.915 -30.765 565.245 -30.435 ;
        RECT 563.555 -30.765 563.885 -30.435 ;
        RECT 558.115 -30.765 558.445 -30.435 ;
        RECT 555.395 -30.765 555.725 -30.435 ;
        RECT 552.675 -30.765 553.005 -30.435 ;
        RECT 551.315 -30.765 551.645 -30.435 ;
        RECT 549.955 -30.765 550.285 -30.435 ;
        RECT 548.595 -30.765 548.925 -30.435 ;
        RECT 543.155 -30.765 543.485 -30.435 ;
        RECT 540.435 -30.765 540.765 -30.435 ;
        RECT 537.715 -30.765 538.045 -30.435 ;
        RECT 536.355 -30.765 536.685 -30.435 ;
        RECT 534.995 -30.765 535.325 -30.435 ;
        RECT 533.635 -30.765 533.965 -30.435 ;
        RECT 528.195 -30.765 528.525 -30.435 ;
        RECT 525.475 -30.765 525.805 -30.435 ;
        RECT 522.755 -30.765 523.085 -30.435 ;
        RECT 521.395 -30.765 521.725 -30.435 ;
        RECT 520.035 -30.765 520.365 -30.435 ;
        RECT 518.675 -30.765 519.005 -30.435 ;
        RECT 513.235 -30.765 513.565 -30.435 ;
        RECT 510.515 -30.765 510.845 -30.435 ;
        RECT 507.795 -30.765 508.125 -30.435 ;
        RECT 506.435 -30.765 506.765 -30.435 ;
        RECT 505.075 -30.765 505.405 -30.435 ;
        RECT 503.715 -30.765 504.045 -30.435 ;
        RECT 498.275 -30.765 498.605 -30.435 ;
        RECT 495.555 -30.765 495.885 -30.435 ;
        RECT 492.835 -30.765 493.165 -30.435 ;
        RECT 491.475 -30.765 491.805 -30.435 ;
        RECT 490.115 -30.765 490.445 -30.435 ;
        RECT 488.755 -30.765 489.085 -30.435 ;
        RECT 483.315 -30.765 483.645 -30.435 ;
        RECT 480.595 -30.765 480.925 -30.435 ;
        RECT 477.875 -30.765 478.205 -30.435 ;
        RECT 476.515 -30.765 476.845 -30.435 ;
        RECT 475.155 -30.765 475.485 -30.435 ;
        RECT 473.795 -30.765 474.125 -30.435 ;
        RECT 468.355 -30.765 468.685 -30.435 ;
        RECT 465.635 -30.765 465.965 -30.435 ;
        RECT 462.915 -30.765 463.245 -30.435 ;
        RECT 461.555 -30.765 461.885 -30.435 ;
        RECT 460.195 -30.765 460.525 -30.435 ;
        RECT 458.835 -30.765 459.165 -30.435 ;
        RECT 453.395 -30.765 453.725 -30.435 ;
        RECT 450.675 -30.765 451.005 -30.435 ;
        RECT 447.955 -30.765 448.285 -30.435 ;
        RECT 446.595 -30.765 446.925 -30.435 ;
        RECT 445.235 -30.765 445.565 -30.435 ;
        RECT 443.875 -30.765 444.205 -30.435 ;
        RECT 438.435 -30.765 438.765 -30.435 ;
        RECT 435.715 -30.765 436.045 -30.435 ;
        RECT 432.995 -30.765 433.325 -30.435 ;
        RECT 431.635 -30.765 431.965 -30.435 ;
        RECT 430.275 -30.765 430.605 -30.435 ;
        RECT 428.915 -30.765 429.245 -30.435 ;
        RECT 423.475 -30.765 423.805 -30.435 ;
        RECT 420.755 -30.765 421.085 -30.435 ;
        RECT 418.035 -30.765 418.365 -30.435 ;
        RECT 416.675 -30.765 417.005 -30.435 ;
        RECT 415.315 -30.765 415.645 -30.435 ;
        RECT 413.955 -30.765 414.285 -30.435 ;
        RECT 408.515 -30.765 408.845 -30.435 ;
        RECT 405.795 -30.765 406.125 -30.435 ;
        RECT 403.075 -30.765 403.405 -30.435 ;
        RECT 401.715 -30.765 402.045 -30.435 ;
        RECT 400.355 -30.765 400.685 -30.435 ;
        RECT 398.995 -30.765 399.325 -30.435 ;
        RECT 393.555 -30.765 393.885 -30.435 ;
        RECT 390.835 -30.765 391.165 -30.435 ;
        RECT 388.115 -30.765 388.445 -30.435 ;
        RECT 386.755 -30.765 387.085 -30.435 ;
        RECT 385.395 -30.765 385.725 -30.435 ;
        RECT 384.035 -30.765 384.365 -30.435 ;
        RECT 378.595 -30.765 378.925 -30.435 ;
        RECT 375.875 -30.765 376.205 -30.435 ;
        RECT 373.155 -30.765 373.485 -30.435 ;
        RECT 371.795 -30.765 372.125 -30.435 ;
        RECT 370.435 -30.765 370.765 -30.435 ;
        RECT 369.075 -30.765 369.405 -30.435 ;
        RECT 363.635 -30.765 363.965 -30.435 ;
        RECT 360.915 -30.765 361.245 -30.435 ;
        RECT 358.195 -30.765 358.525 -30.435 ;
        RECT 356.835 -30.765 357.165 -30.435 ;
        RECT 355.475 -30.765 355.805 -30.435 ;
        RECT 354.115 -30.765 354.445 -30.435 ;
        RECT 351.395 -30.765 351.725 -30.435 ;
        RECT 348.675 -30.765 349.005 -30.435 ;
        RECT 345.955 -30.765 346.285 -30.435 ;
        RECT 343.235 -30.765 343.565 -30.435 ;
        RECT 341.875 -30.765 342.205 -30.435 ;
        RECT 340.515 -30.765 340.845 -30.435 ;
        RECT 339.155 -30.765 339.485 -30.435 ;
        RECT 336.435 -30.765 336.765 -30.435 ;
        RECT 333.715 -30.765 334.045 -30.435 ;
        RECT 330.995 -30.765 331.325 -30.435 ;
        RECT 328.275 -30.765 328.605 -30.435 ;
        RECT 326.915 -30.765 327.245 -30.435 ;
        RECT 325.555 -30.765 325.885 -30.435 ;
        RECT 321.475 -30.765 321.805 -30.435 ;
        RECT 318.755 -30.765 319.085 -30.435 ;
        RECT 316.035 -30.765 316.365 -30.435 ;
        RECT 313.315 -30.765 313.645 -30.435 ;
        RECT 311.955 -30.765 312.285 -30.435 ;
        RECT 310.595 -30.765 310.925 -30.435 ;
        RECT 306.515 -30.765 306.845 -30.435 ;
        RECT 303.795 -30.765 304.125 -30.435 ;
        RECT 301.075 -30.765 301.405 -30.435 ;
        RECT 298.355 -30.765 298.685 -30.435 ;
        RECT 296.995 -30.765 297.325 -30.435 ;
        RECT 295.635 -30.765 295.965 -30.435 ;
        RECT 291.555 -30.765 291.885 -30.435 ;
        RECT 288.835 -30.765 289.165 -30.435 ;
        RECT 284.755 -30.765 285.085 -30.435 ;
        RECT 283.395 -30.765 283.725 -30.435 ;
        RECT 282.035 -30.765 282.365 -30.435 ;
        RECT 280.675 -30.765 281.005 -30.435 ;
        RECT 276.595 -30.765 276.925 -30.435 ;
        RECT 273.875 -30.765 274.205 -30.435 ;
        RECT 272.515 -30.765 272.845 -30.435 ;
        RECT 269.795 -30.765 270.125 -30.435 ;
        RECT 268.435 -30.765 268.765 -30.435 ;
        RECT 267.075 -30.765 267.405 -30.435 ;
        RECT 265.715 -30.765 266.045 -30.435 ;
        RECT 261.635 -30.765 261.965 -30.435 ;
        RECT 257.555 -30.765 257.885 -30.435 ;
        RECT 254.835 -30.765 255.165 -30.435 ;
        RECT 253.475 -30.765 253.805 -30.435 ;
        RECT 252.115 -30.765 252.445 -30.435 ;
        RECT 250.755 -30.765 251.085 -30.435 ;
        RECT 246.675 -30.765 247.005 -30.435 ;
        RECT 242.595 -30.765 242.925 -30.435 ;
        RECT 239.875 -30.765 240.205 -30.435 ;
        RECT 238.515 -30.765 238.845 -30.435 ;
        RECT 237.155 -30.765 237.485 -30.435 ;
        RECT 235.795 -30.765 236.125 -30.435 ;
        RECT 231.715 -30.765 232.045 -30.435 ;
        RECT 227.635 -30.765 227.965 -30.435 ;
        RECT 224.915 -30.765 225.245 -30.435 ;
        RECT 223.555 -30.765 223.885 -30.435 ;
        RECT 222.195 -30.765 222.525 -30.435 ;
        RECT 220.835 -30.765 221.165 -30.435 ;
        RECT 215.395 -30.765 215.725 -30.435 ;
        RECT 212.675 -30.765 213.005 -30.435 ;
        RECT 209.955 -30.765 210.285 -30.435 ;
        RECT 208.595 -30.765 208.925 -30.435 ;
        RECT 207.235 -30.765 207.565 -30.435 ;
        RECT 205.875 -30.765 206.205 -30.435 ;
        RECT 200.435 -30.765 200.765 -30.435 ;
        RECT 197.715 -30.765 198.045 -30.435 ;
        RECT 194.995 -30.765 195.325 -30.435 ;
        RECT 193.635 -30.765 193.965 -30.435 ;
        RECT 192.275 -30.765 192.605 -30.435 ;
        RECT 190.915 -30.765 191.245 -30.435 ;
        RECT 185.475 -30.765 185.805 -30.435 ;
        RECT 182.755 -30.765 183.085 -30.435 ;
        RECT 180.035 -30.765 180.365 -30.435 ;
        RECT 178.675 -30.765 179.005 -30.435 ;
        RECT 177.315 -30.765 177.645 -30.435 ;
        RECT 175.955 -30.765 176.285 -30.435 ;
        RECT 170.515 -30.765 170.845 -30.435 ;
        RECT 167.795 -30.765 168.125 -30.435 ;
        RECT 165.075 -30.765 165.405 -30.435 ;
        RECT 163.715 -30.765 164.045 -30.435 ;
        RECT 162.355 -30.765 162.685 -30.435 ;
        RECT 160.995 -30.765 161.325 -30.435 ;
        RECT 155.555 -30.765 155.885 -30.435 ;
        RECT 152.835 -30.765 153.165 -30.435 ;
        RECT 150.115 -30.765 150.445 -30.435 ;
        RECT 148.755 -30.765 149.085 -30.435 ;
        RECT 147.395 -30.765 147.725 -30.435 ;
        RECT 146.035 -30.765 146.365 -30.435 ;
        RECT 140.595 -30.765 140.925 -30.435 ;
        RECT 137.875 -30.765 138.205 -30.435 ;
        RECT 135.155 -30.765 135.485 -30.435 ;
        RECT 133.795 -30.765 134.125 -30.435 ;
        RECT 132.435 -30.765 132.765 -30.435 ;
        RECT 131.075 -30.765 131.405 -30.435 ;
        RECT 125.635 -30.765 125.965 -30.435 ;
        RECT 122.915 -30.765 123.245 -30.435 ;
        RECT 120.195 -30.765 120.525 -30.435 ;
        RECT 118.835 -30.765 119.165 -30.435 ;
        RECT 117.475 -30.765 117.805 -30.435 ;
        RECT 116.115 -30.765 116.445 -30.435 ;
        RECT 110.675 -30.765 111.005 -30.435 ;
        RECT 107.955 -30.765 108.285 -30.435 ;
        RECT 105.235 -30.765 105.565 -30.435 ;
        RECT 103.875 -30.765 104.205 -30.435 ;
        RECT 102.515 -30.765 102.845 -30.435 ;
        RECT 101.155 -30.765 101.485 -30.435 ;
        RECT 95.715 -30.765 96.045 -30.435 ;
        RECT 92.995 -30.765 93.325 -30.435 ;
        RECT 90.275 -30.765 90.605 -30.435 ;
        RECT 88.915 -30.765 89.245 -30.435 ;
        RECT 87.555 -30.765 87.885 -30.435 ;
        RECT 86.195 -30.765 86.525 -30.435 ;
        RECT 80.755 -30.765 81.085 -30.435 ;
        RECT 78.035 -30.765 78.365 -30.435 ;
        RECT 75.315 -30.765 75.645 -30.435 ;
        RECT 73.955 -30.765 74.285 -30.435 ;
        RECT 72.595 -30.765 72.925 -30.435 ;
        RECT 71.235 -30.765 71.565 -30.435 ;
        RECT 65.795 -30.765 66.125 -30.435 ;
        RECT 63.075 -30.765 63.405 -30.435 ;
        RECT 60.355 -30.765 60.685 -30.435 ;
        RECT 58.995 -30.765 59.325 -30.435 ;
        RECT 57.635 -30.765 57.965 -30.435 ;
        RECT 56.275 -30.765 56.605 -30.435 ;
        RECT 50.835 -30.765 51.165 -30.435 ;
        RECT 48.115 -30.765 48.445 -30.435 ;
        RECT 45.395 -30.765 45.725 -30.435 ;
        RECT 44.035 -30.765 44.365 -30.435 ;
        RECT 42.675 -30.765 43.005 -30.435 ;
        RECT 41.315 -30.765 41.645 -30.435 ;
        RECT 35.875 -30.765 36.205 -30.435 ;
        RECT 33.155 -30.765 33.485 -30.435 ;
        RECT 30.435 -30.765 30.765 -30.435 ;
        RECT 29.075 -30.765 29.405 -30.435 ;
        RECT 27.715 -30.765 28.045 -30.435 ;
        RECT 26.355 -30.765 26.685 -30.435 ;
        RECT 20.915 -30.765 21.245 -30.435 ;
        RECT 18.195 -30.765 18.525 -30.435 ;
        RECT 15.475 -30.765 15.805 -30.435 ;
        RECT 14.115 -30.765 14.445 -30.435 ;
        RECT 12.755 -30.765 13.085 -30.435 ;
        RECT 11.395 -30.765 11.725 -30.435 ;
        RECT 8.675 -30.765 9.005 -30.435 ;
        RECT 7.315 -30.765 7.645 -30.435 ;
        RECT 5.955 -30.765 6.285 -30.435 ;
        RECT 4.595 -30.765 4.925 -30.435 ;
        RECT 3.235 -30.765 3.565 -30.435 ;
        RECT 1.875 -30.765 2.205 -30.435 ;
        RECT 0.515 -30.765 0.845 -30.435 ;
        RECT -0.845 -30.765 -0.515 -30.435 ;
        RECT -1.52 -30.76 954.88 -30.44 ;
        RECT 953.875 -30.765 954.205 -30.435 ;
        RECT 952.515 -30.765 952.845 -30.435 ;
        RECT 951.155 -30.765 951.485 -30.435 ;
        RECT 949.795 -30.765 950.125 -30.435 ;
        RECT 947.075 -30.765 947.405 -30.435 ;
        RECT 945.715 -30.765 946.045 -30.435 ;
        RECT 944.355 -30.765 944.685 -30.435 ;
        RECT 942.995 -30.765 943.325 -30.435 ;
        RECT 941.635 -30.765 941.965 -30.435 ;
        RECT 940.275 -30.765 940.605 -30.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.88 -23.96 778.08 -23.64 ;
        RECT 775.715 -23.965 776.045 -23.635 ;
        RECT 774.355 -23.965 774.685 -23.635 ;
        RECT 772.995 -23.965 773.325 -23.635 ;
        RECT 771.635 -23.965 771.965 -23.635 ;
        RECT 767.555 -23.965 767.885 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.88 -28.04 778.08 -27.72 ;
        RECT 775.715 -28.045 776.045 -27.715 ;
        RECT 774.355 -28.045 774.685 -27.715 ;
        RECT 772.995 -28.045 773.325 -27.715 ;
        RECT 771.635 -28.045 771.965 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 770.96 -34.84 778.08 -34.52 ;
        RECT 777.075 -34.845 777.405 -34.515 ;
        RECT 775.715 -34.845 776.045 -34.515 ;
        RECT 774.355 -34.845 774.685 -34.515 ;
        RECT 772.995 -34.845 773.325 -34.515 ;
        RECT 771.635 -34.845 771.965 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 770.96 -26.68 781.48 -26.36 ;
        RECT 779.795 -26.685 780.125 -26.355 ;
        RECT 775.715 -26.685 776.045 -26.355 ;
        RECT 774.355 -26.685 774.685 -26.355 ;
        RECT 772.995 -26.685 773.325 -26.355 ;
        RECT 771.635 -26.685 771.965 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 785.92 -29.4 792.36 -29.08 ;
        RECT 790.675 -29.405 791.005 -29.075 ;
        RECT 789.315 -29.405 789.645 -29.075 ;
        RECT 787.955 -29.405 788.285 -29.075 ;
        RECT 786.595 -29.405 786.925 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 781.16 -23.96 793.04 -23.64 ;
        RECT 790.675 -23.965 791.005 -23.635 ;
        RECT 789.315 -23.965 789.645 -23.635 ;
        RECT 787.955 -23.965 788.285 -23.635 ;
        RECT 786.595 -23.965 786.925 -23.635 ;
        RECT 782.515 -23.965 782.845 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 781.84 -28.04 793.04 -27.72 ;
        RECT 790.675 -28.045 791.005 -27.715 ;
        RECT 789.315 -28.045 789.645 -27.715 ;
        RECT 787.955 -28.045 788.285 -27.715 ;
        RECT 786.595 -28.045 786.925 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 785.92 -34.84 793.04 -34.52 ;
        RECT 792.035 -34.845 792.365 -34.515 ;
        RECT 790.675 -34.845 791.005 -34.515 ;
        RECT 789.315 -34.845 789.645 -34.515 ;
        RECT 787.955 -34.845 788.285 -34.515 ;
        RECT 786.595 -34.845 786.925 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 785.92 -26.68 796.44 -26.36 ;
        RECT 794.755 -26.685 795.085 -26.355 ;
        RECT 790.675 -26.685 791.005 -26.355 ;
        RECT 789.315 -26.685 789.645 -26.355 ;
        RECT 787.955 -26.685 788.285 -26.355 ;
        RECT 786.595 -26.685 786.925 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 796.12 -23.96 807.32 -23.64 ;
        RECT 805.635 -23.965 805.965 -23.635 ;
        RECT 804.275 -23.965 804.605 -23.635 ;
        RECT 802.915 -23.965 803.245 -23.635 ;
        RECT 801.555 -23.965 801.885 -23.635 ;
        RECT 797.475 -23.965 797.805 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 796.8 -28.04 807.32 -27.72 ;
        RECT 805.635 -28.045 805.965 -27.715 ;
        RECT 804.275 -28.045 804.605 -27.715 ;
        RECT 802.915 -28.045 803.245 -27.715 ;
        RECT 801.555 -28.045 801.885 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 800.88 -29.4 807.32 -29.08 ;
        RECT 805.635 -29.405 805.965 -29.075 ;
        RECT 804.275 -29.405 804.605 -29.075 ;
        RECT 802.915 -29.405 803.245 -29.075 ;
        RECT 801.555 -29.405 801.885 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 806.995 -34.845 807.325 -34.515 ;
        RECT 800.88 -34.84 807.325 -34.52 ;
        RECT 805.635 -34.845 805.965 -34.515 ;
        RECT 804.275 -34.845 804.605 -34.515 ;
        RECT 802.915 -34.845 803.245 -34.515 ;
        RECT 801.555 -34.845 801.885 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 800.88 -26.68 811.4 -26.36 ;
        RECT 809.715 -26.685 810.045 -26.355 ;
        RECT 805.635 -26.685 805.965 -26.355 ;
        RECT 804.275 -26.685 804.605 -26.355 ;
        RECT 802.915 -26.685 803.245 -26.355 ;
        RECT 801.555 -26.685 801.885 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 815.84 -29.4 821.6 -29.08 ;
        RECT 820.595 -29.405 820.925 -29.075 ;
        RECT 819.235 -29.405 819.565 -29.075 ;
        RECT 817.875 -29.405 818.205 -29.075 ;
        RECT 816.515 -29.405 816.845 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 811.08 -23.96 822.28 -23.64 ;
        RECT 820.595 -23.965 820.925 -23.635 ;
        RECT 819.235 -23.965 819.565 -23.635 ;
        RECT 817.875 -23.965 818.205 -23.635 ;
        RECT 816.515 -23.965 816.845 -23.635 ;
        RECT 812.435 -23.965 812.765 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 811.76 -28.04 822.28 -27.72 ;
        RECT 820.595 -28.045 820.925 -27.715 ;
        RECT 819.235 -28.045 819.565 -27.715 ;
        RECT 817.875 -28.045 818.205 -27.715 ;
        RECT 816.515 -28.045 816.845 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 821.955 -34.845 822.285 -34.515 ;
        RECT 815.84 -34.84 822.285 -34.52 ;
        RECT 820.595 -34.845 820.925 -34.515 ;
        RECT 819.235 -34.845 819.565 -34.515 ;
        RECT 817.875 -34.845 818.205 -34.515 ;
        RECT 816.515 -34.845 816.845 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 815.84 -26.68 826.36 -26.36 ;
        RECT 824.675 -26.685 825.005 -26.355 ;
        RECT 823.315 -26.685 823.645 -26.355 ;
        RECT 820.595 -26.685 820.925 -26.355 ;
        RECT 819.235 -26.685 819.565 -26.355 ;
        RECT 817.875 -26.685 818.205 -26.355 ;
        RECT 816.515 -26.685 816.845 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 830.8 -29.4 836.56 -29.08 ;
        RECT 835.555 -29.405 835.885 -29.075 ;
        RECT 834.195 -29.405 834.525 -29.075 ;
        RECT 832.835 -29.405 833.165 -29.075 ;
        RECT 831.475 -29.405 831.805 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 826.04 -23.96 837.24 -23.64 ;
        RECT 835.555 -23.965 835.885 -23.635 ;
        RECT 834.195 -23.965 834.525 -23.635 ;
        RECT 832.835 -23.965 833.165 -23.635 ;
        RECT 831.475 -23.965 831.805 -23.635 ;
        RECT 827.395 -23.965 827.725 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 826.72 -28.04 837.24 -27.72 ;
        RECT 835.555 -28.045 835.885 -27.715 ;
        RECT 834.195 -28.045 834.525 -27.715 ;
        RECT 832.835 -28.045 833.165 -27.715 ;
        RECT 831.475 -28.045 831.805 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 836.915 -34.845 837.245 -34.515 ;
        RECT 830.8 -34.84 837.245 -34.52 ;
        RECT 835.555 -34.845 835.885 -34.515 ;
        RECT 834.195 -34.845 834.525 -34.515 ;
        RECT 832.835 -34.845 833.165 -34.515 ;
        RECT 831.475 -34.845 831.805 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 830.8 -26.68 841.32 -26.36 ;
        RECT 839.635 -26.685 839.965 -26.355 ;
        RECT 838.275 -26.685 838.605 -26.355 ;
        RECT 835.555 -26.685 835.885 -26.355 ;
        RECT 834.195 -26.685 834.525 -26.355 ;
        RECT 832.835 -26.685 833.165 -26.355 ;
        RECT 831.475 -26.685 831.805 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 845.76 -29.4 851.52 -29.08 ;
        RECT 850.515 -29.405 850.845 -29.075 ;
        RECT 849.155 -29.405 849.485 -29.075 ;
        RECT 847.795 -29.405 848.125 -29.075 ;
        RECT 846.435 -29.405 846.765 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 841 -23.96 852.2 -23.64 ;
        RECT 850.515 -23.965 850.845 -23.635 ;
        RECT 849.155 -23.965 849.485 -23.635 ;
        RECT 847.795 -23.965 848.125 -23.635 ;
        RECT 846.435 -23.965 846.765 -23.635 ;
        RECT 842.355 -23.965 842.685 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 841.68 -28.04 852.2 -27.72 ;
        RECT 850.515 -28.045 850.845 -27.715 ;
        RECT 849.155 -28.045 849.485 -27.715 ;
        RECT 847.795 -28.045 848.125 -27.715 ;
        RECT 846.435 -28.045 846.765 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 851.875 -34.845 852.205 -34.515 ;
        RECT 845.76 -34.84 852.205 -34.52 ;
        RECT 850.515 -34.845 850.845 -34.515 ;
        RECT 849.155 -34.845 849.485 -34.515 ;
        RECT 847.795 -34.845 848.125 -34.515 ;
        RECT 846.435 -34.845 846.765 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 845.76 -26.68 856.28 -26.36 ;
        RECT 854.595 -26.685 854.925 -26.355 ;
        RECT 853.235 -26.685 853.565 -26.355 ;
        RECT 850.515 -26.685 850.845 -26.355 ;
        RECT 849.155 -26.685 849.485 -26.355 ;
        RECT 847.795 -26.685 848.125 -26.355 ;
        RECT 846.435 -26.685 846.765 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 860.04 -29.4 866.48 -29.08 ;
        RECT 865.475 -29.405 865.805 -29.075 ;
        RECT 864.115 -29.405 864.445 -29.075 ;
        RECT 862.755 -29.405 863.085 -29.075 ;
        RECT 861.395 -29.405 861.725 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 855.96 -23.96 867.16 -23.64 ;
        RECT 865.475 -23.965 865.805 -23.635 ;
        RECT 864.115 -23.965 864.445 -23.635 ;
        RECT 862.755 -23.965 863.085 -23.635 ;
        RECT 861.395 -23.965 861.725 -23.635 ;
        RECT 860.035 -23.965 860.365 -23.635 ;
        RECT 857.315 -23.965 857.645 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 856.64 -28.04 867.16 -27.72 ;
        RECT 865.475 -28.045 865.805 -27.715 ;
        RECT 864.115 -28.045 864.445 -27.715 ;
        RECT 862.755 -28.045 863.085 -27.715 ;
        RECT 861.395 -28.045 861.725 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 866.835 -34.845 867.165 -34.515 ;
        RECT 860.04 -34.84 867.165 -34.52 ;
        RECT 865.475 -34.845 865.805 -34.515 ;
        RECT 864.115 -34.845 864.445 -34.515 ;
        RECT 862.755 -34.845 863.085 -34.515 ;
        RECT 861.395 -34.845 861.725 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 860.04 -26.68 871.24 -26.36 ;
        RECT 869.555 -26.685 869.885 -26.355 ;
        RECT 868.195 -26.685 868.525 -26.355 ;
        RECT 865.475 -26.685 865.805 -26.355 ;
        RECT 864.115 -26.685 864.445 -26.355 ;
        RECT 862.755 -26.685 863.085 -26.355 ;
        RECT 861.395 -26.685 861.725 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 875 -29.4 881.44 -29.08 ;
        RECT 880.435 -29.405 880.765 -29.075 ;
        RECT 879.075 -29.405 879.405 -29.075 ;
        RECT 877.715 -29.405 878.045 -29.075 ;
        RECT 876.355 -29.405 876.685 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 870.92 -23.96 882.12 -23.64 ;
        RECT 880.435 -23.965 880.765 -23.635 ;
        RECT 879.075 -23.965 879.405 -23.635 ;
        RECT 877.715 -23.965 878.045 -23.635 ;
        RECT 876.355 -23.965 876.685 -23.635 ;
        RECT 874.995 -23.965 875.325 -23.635 ;
        RECT 872.275 -23.965 872.605 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 871.6 -28.04 882.12 -27.72 ;
        RECT 880.435 -28.045 880.765 -27.715 ;
        RECT 879.075 -28.045 879.405 -27.715 ;
        RECT 877.715 -28.045 878.045 -27.715 ;
        RECT 876.355 -28.045 876.685 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 881.795 -34.845 882.125 -34.515 ;
        RECT 875 -34.84 882.125 -34.52 ;
        RECT 880.435 -34.845 880.765 -34.515 ;
        RECT 879.075 -34.845 879.405 -34.515 ;
        RECT 877.715 -34.845 878.045 -34.515 ;
        RECT 876.355 -34.845 876.685 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 875 -26.68 886.2 -26.36 ;
        RECT 884.515 -26.685 884.845 -26.355 ;
        RECT 883.155 -26.685 883.485 -26.355 ;
        RECT 880.435 -26.685 880.765 -26.355 ;
        RECT 879.075 -26.685 879.405 -26.355 ;
        RECT 877.715 -26.685 878.045 -26.355 ;
        RECT 876.355 -26.685 876.685 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 889.96 -29.4 896.4 -29.08 ;
        RECT 895.395 -29.405 895.725 -29.075 ;
        RECT 894.035 -29.405 894.365 -29.075 ;
        RECT 892.675 -29.405 893.005 -29.075 ;
        RECT 891.315 -29.405 891.645 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 885.88 -23.96 897.08 -23.64 ;
        RECT 895.395 -23.965 895.725 -23.635 ;
        RECT 894.035 -23.965 894.365 -23.635 ;
        RECT 892.675 -23.965 893.005 -23.635 ;
        RECT 891.315 -23.965 891.645 -23.635 ;
        RECT 889.955 -23.965 890.285 -23.635 ;
        RECT 887.235 -23.965 887.565 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 886.56 -28.04 897.08 -27.72 ;
        RECT 895.395 -28.045 895.725 -27.715 ;
        RECT 894.035 -28.045 894.365 -27.715 ;
        RECT 892.675 -28.045 893.005 -27.715 ;
        RECT 891.315 -28.045 891.645 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 896.755 -34.845 897.085 -34.515 ;
        RECT 889.96 -34.84 897.085 -34.52 ;
        RECT 895.395 -34.845 895.725 -34.515 ;
        RECT 894.035 -34.845 894.365 -34.515 ;
        RECT 892.675 -34.845 893.005 -34.515 ;
        RECT 891.315 -34.845 891.645 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 889.96 -26.68 900.48 -26.36 ;
        RECT 899.475 -26.685 899.805 -26.355 ;
        RECT 898.115 -26.685 898.445 -26.355 ;
        RECT 895.395 -26.685 895.725 -26.355 ;
        RECT 894.035 -26.685 894.365 -26.355 ;
        RECT 892.675 -26.685 893.005 -26.355 ;
        RECT 891.315 -26.685 891.645 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 904.92 -29.4 911.36 -29.08 ;
        RECT 910.355 -29.405 910.685 -29.075 ;
        RECT 908.995 -29.405 909.325 -29.075 ;
        RECT 907.635 -29.405 907.965 -29.075 ;
        RECT 906.275 -29.405 906.605 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 900.84 -23.96 912.04 -23.64 ;
        RECT 910.355 -23.965 910.685 -23.635 ;
        RECT 908.995 -23.965 909.325 -23.635 ;
        RECT 907.635 -23.965 907.965 -23.635 ;
        RECT 906.275 -23.965 906.605 -23.635 ;
        RECT 904.915 -23.965 905.245 -23.635 ;
        RECT 902.195 -23.965 902.525 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 901.52 -28.04 912.04 -27.72 ;
        RECT 910.355 -28.045 910.685 -27.715 ;
        RECT 908.995 -28.045 909.325 -27.715 ;
        RECT 907.635 -28.045 907.965 -27.715 ;
        RECT 906.275 -28.045 906.605 -27.715 ;
        RECT 902.195 -28.045 902.525 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 911.715 -34.845 912.045 -34.515 ;
        RECT 904.92 -34.84 912.045 -34.52 ;
        RECT 910.355 -34.845 910.685 -34.515 ;
        RECT 908.995 -34.845 909.325 -34.515 ;
        RECT 907.635 -34.845 907.965 -34.515 ;
        RECT 906.275 -34.845 906.605 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 904.92 -26.68 915.44 -26.36 ;
        RECT 914.435 -26.685 914.765 -26.355 ;
        RECT 913.075 -26.685 913.405 -26.355 ;
        RECT 910.355 -26.685 910.685 -26.355 ;
        RECT 908.995 -26.685 909.325 -26.355 ;
        RECT 907.635 -26.685 907.965 -26.355 ;
        RECT 906.275 -26.685 906.605 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 923.955 -19.885 924.285 -19.555 ;
        RECT -1.52 -19.88 924.285 -19.56 ;
        RECT 922.595 -19.885 922.925 -19.555 ;
        RECT 921.235 -19.885 921.565 -19.555 ;
        RECT 919.875 -19.885 920.205 -19.555 ;
        RECT 918.515 -19.885 918.845 -19.555 ;
        RECT 917.155 -19.885 917.485 -19.555 ;
        RECT 913.075 -19.885 913.405 -19.555 ;
        RECT 910.355 -19.885 910.685 -19.555 ;
        RECT 908.995 -19.885 909.325 -19.555 ;
        RECT 907.635 -19.885 907.965 -19.555 ;
        RECT 906.275 -19.885 906.605 -19.555 ;
        RECT 904.915 -19.885 905.245 -19.555 ;
        RECT 903.555 -19.885 903.885 -19.555 ;
        RECT 902.195 -19.885 902.525 -19.555 ;
        RECT 898.115 -19.885 898.445 -19.555 ;
        RECT 895.395 -19.885 895.725 -19.555 ;
        RECT 894.035 -19.885 894.365 -19.555 ;
        RECT 892.675 -19.885 893.005 -19.555 ;
        RECT 891.315 -19.885 891.645 -19.555 ;
        RECT 889.955 -19.885 890.285 -19.555 ;
        RECT 888.595 -19.885 888.925 -19.555 ;
        RECT 887.235 -19.885 887.565 -19.555 ;
        RECT 883.155 -19.885 883.485 -19.555 ;
        RECT 880.435 -19.885 880.765 -19.555 ;
        RECT 879.075 -19.885 879.405 -19.555 ;
        RECT 877.715 -19.885 878.045 -19.555 ;
        RECT 876.355 -19.885 876.685 -19.555 ;
        RECT 874.995 -19.885 875.325 -19.555 ;
        RECT 873.635 -19.885 873.965 -19.555 ;
        RECT 872.275 -19.885 872.605 -19.555 ;
        RECT 868.195 -19.885 868.525 -19.555 ;
        RECT 865.475 -19.885 865.805 -19.555 ;
        RECT 864.115 -19.885 864.445 -19.555 ;
        RECT 862.755 -19.885 863.085 -19.555 ;
        RECT 861.395 -19.885 861.725 -19.555 ;
        RECT 860.035 -19.885 860.365 -19.555 ;
        RECT 858.675 -19.885 859.005 -19.555 ;
        RECT 857.315 -19.885 857.645 -19.555 ;
        RECT 853.235 -19.885 853.565 -19.555 ;
        RECT 850.515 -19.885 850.845 -19.555 ;
        RECT 849.155 -19.885 849.485 -19.555 ;
        RECT 847.795 -19.885 848.125 -19.555 ;
        RECT 846.435 -19.885 846.765 -19.555 ;
        RECT 845.075 -19.885 845.405 -19.555 ;
        RECT 843.715 -19.885 844.045 -19.555 ;
        RECT 842.355 -19.885 842.685 -19.555 ;
        RECT 838.275 -19.885 838.605 -19.555 ;
        RECT 835.555 -19.885 835.885 -19.555 ;
        RECT 834.195 -19.885 834.525 -19.555 ;
        RECT 832.835 -19.885 833.165 -19.555 ;
        RECT 831.475 -19.885 831.805 -19.555 ;
        RECT 830.115 -19.885 830.445 -19.555 ;
        RECT 828.755 -19.885 829.085 -19.555 ;
        RECT 827.395 -19.885 827.725 -19.555 ;
        RECT 823.315 -19.885 823.645 -19.555 ;
        RECT 820.595 -19.885 820.925 -19.555 ;
        RECT 819.235 -19.885 819.565 -19.555 ;
        RECT 817.875 -19.885 818.205 -19.555 ;
        RECT 816.515 -19.885 816.845 -19.555 ;
        RECT 815.155 -19.885 815.485 -19.555 ;
        RECT 813.795 -19.885 814.125 -19.555 ;
        RECT 812.435 -19.885 812.765 -19.555 ;
        RECT 806.995 -19.885 807.325 -19.555 ;
        RECT 805.635 -19.885 805.965 -19.555 ;
        RECT 804.275 -19.885 804.605 -19.555 ;
        RECT 802.915 -19.885 803.245 -19.555 ;
        RECT 801.555 -19.885 801.885 -19.555 ;
        RECT 800.195 -19.885 800.525 -19.555 ;
        RECT 798.835 -19.885 799.165 -19.555 ;
        RECT 797.475 -19.885 797.805 -19.555 ;
        RECT 792.035 -19.885 792.365 -19.555 ;
        RECT 790.675 -19.885 791.005 -19.555 ;
        RECT 789.315 -19.885 789.645 -19.555 ;
        RECT 787.955 -19.885 788.285 -19.555 ;
        RECT 786.595 -19.885 786.925 -19.555 ;
        RECT 785.235 -19.885 785.565 -19.555 ;
        RECT 783.875 -19.885 784.205 -19.555 ;
        RECT 782.515 -19.885 782.845 -19.555 ;
        RECT 777.075 -19.885 777.405 -19.555 ;
        RECT 775.715 -19.885 776.045 -19.555 ;
        RECT 774.355 -19.885 774.685 -19.555 ;
        RECT 772.995 -19.885 773.325 -19.555 ;
        RECT 771.635 -19.885 771.965 -19.555 ;
        RECT 770.275 -19.885 770.605 -19.555 ;
        RECT 768.915 -19.885 769.245 -19.555 ;
        RECT 767.555 -19.885 767.885 -19.555 ;
        RECT 762.115 -19.885 762.445 -19.555 ;
        RECT 760.755 -19.885 761.085 -19.555 ;
        RECT 759.395 -19.885 759.725 -19.555 ;
        RECT 758.035 -19.885 758.365 -19.555 ;
        RECT 756.675 -19.885 757.005 -19.555 ;
        RECT 755.315 -19.885 755.645 -19.555 ;
        RECT 753.955 -19.885 754.285 -19.555 ;
        RECT 752.595 -19.885 752.925 -19.555 ;
        RECT 747.155 -19.885 747.485 -19.555 ;
        RECT 745.795 -19.885 746.125 -19.555 ;
        RECT 744.435 -19.885 744.765 -19.555 ;
        RECT 743.075 -19.885 743.405 -19.555 ;
        RECT 741.715 -19.885 742.045 -19.555 ;
        RECT 740.355 -19.885 740.685 -19.555 ;
        RECT 738.995 -19.885 739.325 -19.555 ;
        RECT 737.635 -19.885 737.965 -19.555 ;
        RECT 732.195 -19.885 732.525 -19.555 ;
        RECT 730.835 -19.885 731.165 -19.555 ;
        RECT 729.475 -19.885 729.805 -19.555 ;
        RECT 728.115 -19.885 728.445 -19.555 ;
        RECT 726.755 -19.885 727.085 -19.555 ;
        RECT 725.395 -19.885 725.725 -19.555 ;
        RECT 724.035 -19.885 724.365 -19.555 ;
        RECT 722.675 -19.885 723.005 -19.555 ;
        RECT 717.235 -19.885 717.565 -19.555 ;
        RECT 715.875 -19.885 716.205 -19.555 ;
        RECT 714.515 -19.885 714.845 -19.555 ;
        RECT 713.155 -19.885 713.485 -19.555 ;
        RECT 711.795 -19.885 712.125 -19.555 ;
        RECT 710.435 -19.885 710.765 -19.555 ;
        RECT 709.075 -19.885 709.405 -19.555 ;
        RECT 707.715 -19.885 708.045 -19.555 ;
        RECT 702.275 -19.885 702.605 -19.555 ;
        RECT 700.915 -19.885 701.245 -19.555 ;
        RECT 699.555 -19.885 699.885 -19.555 ;
        RECT 698.195 -19.885 698.525 -19.555 ;
        RECT 696.835 -19.885 697.165 -19.555 ;
        RECT 695.475 -19.885 695.805 -19.555 ;
        RECT 694.115 -19.885 694.445 -19.555 ;
        RECT 692.755 -19.885 693.085 -19.555 ;
        RECT 687.315 -19.885 687.645 -19.555 ;
        RECT 685.955 -19.885 686.285 -19.555 ;
        RECT 684.595 -19.885 684.925 -19.555 ;
        RECT 683.235 -19.885 683.565 -19.555 ;
        RECT 681.875 -19.885 682.205 -19.555 ;
        RECT 680.515 -19.885 680.845 -19.555 ;
        RECT 679.155 -19.885 679.485 -19.555 ;
        RECT 677.795 -19.885 678.125 -19.555 ;
        RECT 672.355 -19.885 672.685 -19.555 ;
        RECT 670.995 -19.885 671.325 -19.555 ;
        RECT 669.635 -19.885 669.965 -19.555 ;
        RECT 668.275 -19.885 668.605 -19.555 ;
        RECT 666.915 -19.885 667.245 -19.555 ;
        RECT 665.555 -19.885 665.885 -19.555 ;
        RECT 664.195 -19.885 664.525 -19.555 ;
        RECT 662.835 -19.885 663.165 -19.555 ;
        RECT 657.395 -19.885 657.725 -19.555 ;
        RECT 656.035 -19.885 656.365 -19.555 ;
        RECT 654.675 -19.885 655.005 -19.555 ;
        RECT 653.315 -19.885 653.645 -19.555 ;
        RECT 651.955 -19.885 652.285 -19.555 ;
        RECT 650.595 -19.885 650.925 -19.555 ;
        RECT 649.235 -19.885 649.565 -19.555 ;
        RECT 647.875 -19.885 648.205 -19.555 ;
        RECT 642.435 -19.885 642.765 -19.555 ;
        RECT 641.075 -19.885 641.405 -19.555 ;
        RECT 639.715 -19.885 640.045 -19.555 ;
        RECT 638.355 -19.885 638.685 -19.555 ;
        RECT 636.995 -19.885 637.325 -19.555 ;
        RECT 635.635 -19.885 635.965 -19.555 ;
        RECT 634.275 -19.885 634.605 -19.555 ;
        RECT 632.915 -19.885 633.245 -19.555 ;
        RECT 627.475 -19.885 627.805 -19.555 ;
        RECT 626.115 -19.885 626.445 -19.555 ;
        RECT 624.755 -19.885 625.085 -19.555 ;
        RECT 623.395 -19.885 623.725 -19.555 ;
        RECT 622.035 -19.885 622.365 -19.555 ;
        RECT 620.675 -19.885 621.005 -19.555 ;
        RECT 619.315 -19.885 619.645 -19.555 ;
        RECT 617.955 -19.885 618.285 -19.555 ;
        RECT 612.515 -19.885 612.845 -19.555 ;
        RECT 611.155 -19.885 611.485 -19.555 ;
        RECT 609.795 -19.885 610.125 -19.555 ;
        RECT 608.435 -19.885 608.765 -19.555 ;
        RECT 607.075 -19.885 607.405 -19.555 ;
        RECT 605.715 -19.885 606.045 -19.555 ;
        RECT 604.355 -19.885 604.685 -19.555 ;
        RECT 602.995 -19.885 603.325 -19.555 ;
        RECT 600.275 -19.885 600.605 -19.555 ;
        RECT 597.555 -19.885 597.885 -19.555 ;
        RECT 596.195 -19.885 596.525 -19.555 ;
        RECT 594.835 -19.885 595.165 -19.555 ;
        RECT 593.475 -19.885 593.805 -19.555 ;
        RECT 592.115 -19.885 592.445 -19.555 ;
        RECT 590.755 -19.885 591.085 -19.555 ;
        RECT 589.395 -19.885 589.725 -19.555 ;
        RECT 588.035 -19.885 588.365 -19.555 ;
        RECT 585.315 -19.885 585.645 -19.555 ;
        RECT 582.595 -19.885 582.925 -19.555 ;
        RECT 581.235 -19.885 581.565 -19.555 ;
        RECT 579.875 -19.885 580.205 -19.555 ;
        RECT 578.515 -19.885 578.845 -19.555 ;
        RECT 577.155 -19.885 577.485 -19.555 ;
        RECT 575.795 -19.885 576.125 -19.555 ;
        RECT 574.435 -19.885 574.765 -19.555 ;
        RECT 570.355 -19.885 570.685 -19.555 ;
        RECT 567.635 -19.885 567.965 -19.555 ;
        RECT 566.275 -19.885 566.605 -19.555 ;
        RECT 564.915 -19.885 565.245 -19.555 ;
        RECT 563.555 -19.885 563.885 -19.555 ;
        RECT 562.195 -19.885 562.525 -19.555 ;
        RECT 560.835 -19.885 561.165 -19.555 ;
        RECT 559.475 -19.885 559.805 -19.555 ;
        RECT 555.395 -19.885 555.725 -19.555 ;
        RECT 552.675 -19.885 553.005 -19.555 ;
        RECT 551.315 -19.885 551.645 -19.555 ;
        RECT 549.955 -19.885 550.285 -19.555 ;
        RECT 548.595 -19.885 548.925 -19.555 ;
        RECT 547.235 -19.885 547.565 -19.555 ;
        RECT 545.875 -19.885 546.205 -19.555 ;
        RECT 544.515 -19.885 544.845 -19.555 ;
        RECT 540.435 -19.885 540.765 -19.555 ;
        RECT 537.715 -19.885 538.045 -19.555 ;
        RECT 536.355 -19.885 536.685 -19.555 ;
        RECT 534.995 -19.885 535.325 -19.555 ;
        RECT 533.635 -19.885 533.965 -19.555 ;
        RECT 532.275 -19.885 532.605 -19.555 ;
        RECT 530.915 -19.885 531.245 -19.555 ;
        RECT 529.555 -19.885 529.885 -19.555 ;
        RECT 525.475 -19.885 525.805 -19.555 ;
        RECT 522.755 -19.885 523.085 -19.555 ;
        RECT 521.395 -19.885 521.725 -19.555 ;
        RECT 520.035 -19.885 520.365 -19.555 ;
        RECT 518.675 -19.885 519.005 -19.555 ;
        RECT 517.315 -19.885 517.645 -19.555 ;
        RECT 515.955 -19.885 516.285 -19.555 ;
        RECT 514.595 -19.885 514.925 -19.555 ;
        RECT 510.515 -19.885 510.845 -19.555 ;
        RECT 507.795 -19.885 508.125 -19.555 ;
        RECT 506.435 -19.885 506.765 -19.555 ;
        RECT 505.075 -19.885 505.405 -19.555 ;
        RECT 503.715 -19.885 504.045 -19.555 ;
        RECT 502.355 -19.885 502.685 -19.555 ;
        RECT 500.995 -19.885 501.325 -19.555 ;
        RECT 499.635 -19.885 499.965 -19.555 ;
        RECT 495.555 -19.885 495.885 -19.555 ;
        RECT 492.835 -19.885 493.165 -19.555 ;
        RECT 491.475 -19.885 491.805 -19.555 ;
        RECT 490.115 -19.885 490.445 -19.555 ;
        RECT 488.755 -19.885 489.085 -19.555 ;
        RECT 487.395 -19.885 487.725 -19.555 ;
        RECT 486.035 -19.885 486.365 -19.555 ;
        RECT 484.675 -19.885 485.005 -19.555 ;
        RECT 480.595 -19.885 480.925 -19.555 ;
        RECT 477.875 -19.885 478.205 -19.555 ;
        RECT 476.515 -19.885 476.845 -19.555 ;
        RECT 475.155 -19.885 475.485 -19.555 ;
        RECT 473.795 -19.885 474.125 -19.555 ;
        RECT 472.435 -19.885 472.765 -19.555 ;
        RECT 471.075 -19.885 471.405 -19.555 ;
        RECT 469.715 -19.885 470.045 -19.555 ;
        RECT 464.275 -19.885 464.605 -19.555 ;
        RECT 462.915 -19.885 463.245 -19.555 ;
        RECT 461.555 -19.885 461.885 -19.555 ;
        RECT 460.195 -19.885 460.525 -19.555 ;
        RECT 458.835 -19.885 459.165 -19.555 ;
        RECT 457.475 -19.885 457.805 -19.555 ;
        RECT 456.115 -19.885 456.445 -19.555 ;
        RECT 454.755 -19.885 455.085 -19.555 ;
        RECT 449.315 -19.885 449.645 -19.555 ;
        RECT 447.955 -19.885 448.285 -19.555 ;
        RECT 446.595 -19.885 446.925 -19.555 ;
        RECT 445.235 -19.885 445.565 -19.555 ;
        RECT 443.875 -19.885 444.205 -19.555 ;
        RECT 442.515 -19.885 442.845 -19.555 ;
        RECT 441.155 -19.885 441.485 -19.555 ;
        RECT 439.795 -19.885 440.125 -19.555 ;
        RECT 434.355 -19.885 434.685 -19.555 ;
        RECT 432.995 -19.885 433.325 -19.555 ;
        RECT 431.635 -19.885 431.965 -19.555 ;
        RECT 430.275 -19.885 430.605 -19.555 ;
        RECT 428.915 -19.885 429.245 -19.555 ;
        RECT 427.555 -19.885 427.885 -19.555 ;
        RECT 426.195 -19.885 426.525 -19.555 ;
        RECT 424.835 -19.885 425.165 -19.555 ;
        RECT 419.395 -19.885 419.725 -19.555 ;
        RECT 418.035 -19.885 418.365 -19.555 ;
        RECT 416.675 -19.885 417.005 -19.555 ;
        RECT 415.315 -19.885 415.645 -19.555 ;
        RECT 413.955 -19.885 414.285 -19.555 ;
        RECT 412.595 -19.885 412.925 -19.555 ;
        RECT 411.235 -19.885 411.565 -19.555 ;
        RECT 409.875 -19.885 410.205 -19.555 ;
        RECT 404.435 -19.885 404.765 -19.555 ;
        RECT 403.075 -19.885 403.405 -19.555 ;
        RECT 401.715 -19.885 402.045 -19.555 ;
        RECT 400.355 -19.885 400.685 -19.555 ;
        RECT 398.995 -19.885 399.325 -19.555 ;
        RECT 397.635 -19.885 397.965 -19.555 ;
        RECT 396.275 -19.885 396.605 -19.555 ;
        RECT 394.915 -19.885 395.245 -19.555 ;
        RECT 389.475 -19.885 389.805 -19.555 ;
        RECT 388.115 -19.885 388.445 -19.555 ;
        RECT 386.755 -19.885 387.085 -19.555 ;
        RECT 385.395 -19.885 385.725 -19.555 ;
        RECT 384.035 -19.885 384.365 -19.555 ;
        RECT 382.675 -19.885 383.005 -19.555 ;
        RECT 381.315 -19.885 381.645 -19.555 ;
        RECT 379.955 -19.885 380.285 -19.555 ;
        RECT 374.515 -19.885 374.845 -19.555 ;
        RECT 373.155 -19.885 373.485 -19.555 ;
        RECT 371.795 -19.885 372.125 -19.555 ;
        RECT 370.435 -19.885 370.765 -19.555 ;
        RECT 369.075 -19.885 369.405 -19.555 ;
        RECT 367.715 -19.885 368.045 -19.555 ;
        RECT 366.355 -19.885 366.685 -19.555 ;
        RECT 364.995 -19.885 365.325 -19.555 ;
        RECT 359.555 -19.885 359.885 -19.555 ;
        RECT 358.195 -19.885 358.525 -19.555 ;
        RECT 356.835 -19.885 357.165 -19.555 ;
        RECT 355.475 -19.885 355.805 -19.555 ;
        RECT 354.115 -19.885 354.445 -19.555 ;
        RECT 352.755 -19.885 353.085 -19.555 ;
        RECT 351.395 -19.885 351.725 -19.555 ;
        RECT 350.035 -19.885 350.365 -19.555 ;
        RECT 344.595 -19.885 344.925 -19.555 ;
        RECT 343.235 -19.885 343.565 -19.555 ;
        RECT 341.875 -19.885 342.205 -19.555 ;
        RECT 340.515 -19.885 340.845 -19.555 ;
        RECT 339.155 -19.885 339.485 -19.555 ;
        RECT 337.795 -19.885 338.125 -19.555 ;
        RECT 336.435 -19.885 336.765 -19.555 ;
        RECT 335.075 -19.885 335.405 -19.555 ;
        RECT 329.635 -19.885 329.965 -19.555 ;
        RECT 328.275 -19.885 328.605 -19.555 ;
        RECT 326.915 -19.885 327.245 -19.555 ;
        RECT 325.555 -19.885 325.885 -19.555 ;
        RECT 324.195 -19.885 324.525 -19.555 ;
        RECT 322.835 -19.885 323.165 -19.555 ;
        RECT 321.475 -19.885 321.805 -19.555 ;
        RECT 320.115 -19.885 320.445 -19.555 ;
        RECT 314.675 -19.885 315.005 -19.555 ;
        RECT 313.315 -19.885 313.645 -19.555 ;
        RECT 311.955 -19.885 312.285 -19.555 ;
        RECT 310.595 -19.885 310.925 -19.555 ;
        RECT 309.235 -19.885 309.565 -19.555 ;
        RECT 307.875 -19.885 308.205 -19.555 ;
        RECT 306.515 -19.885 306.845 -19.555 ;
        RECT 305.155 -19.885 305.485 -19.555 ;
        RECT 299.715 -19.885 300.045 -19.555 ;
        RECT 298.355 -19.885 298.685 -19.555 ;
        RECT 296.995 -19.885 297.325 -19.555 ;
        RECT 295.635 -19.885 295.965 -19.555 ;
        RECT 294.275 -19.885 294.605 -19.555 ;
        RECT 292.915 -19.885 293.245 -19.555 ;
        RECT 291.555 -19.885 291.885 -19.555 ;
        RECT 290.195 -19.885 290.525 -19.555 ;
        RECT 284.755 -19.885 285.085 -19.555 ;
        RECT 283.395 -19.885 283.725 -19.555 ;
        RECT 282.035 -19.885 282.365 -19.555 ;
        RECT 280.675 -19.885 281.005 -19.555 ;
        RECT 279.315 -19.885 279.645 -19.555 ;
        RECT 277.955 -19.885 278.285 -19.555 ;
        RECT 276.595 -19.885 276.925 -19.555 ;
        RECT 275.235 -19.885 275.565 -19.555 ;
        RECT 272.515 -19.885 272.845 -19.555 ;
        RECT 269.795 -19.885 270.125 -19.555 ;
        RECT 268.435 -19.885 268.765 -19.555 ;
        RECT 267.075 -19.885 267.405 -19.555 ;
        RECT 265.715 -19.885 266.045 -19.555 ;
        RECT 264.355 -19.885 264.685 -19.555 ;
        RECT 262.995 -19.885 263.325 -19.555 ;
        RECT 261.635 -19.885 261.965 -19.555 ;
        RECT 260.275 -19.885 260.605 -19.555 ;
        RECT 257.555 -19.885 257.885 -19.555 ;
        RECT 254.835 -19.885 255.165 -19.555 ;
        RECT 253.475 -19.885 253.805 -19.555 ;
        RECT 252.115 -19.885 252.445 -19.555 ;
        RECT 250.755 -19.885 251.085 -19.555 ;
        RECT 249.395 -19.885 249.725 -19.555 ;
        RECT 248.035 -19.885 248.365 -19.555 ;
        RECT 246.675 -19.885 247.005 -19.555 ;
        RECT 242.595 -19.885 242.925 -19.555 ;
        RECT 239.875 -19.885 240.205 -19.555 ;
        RECT 238.515 -19.885 238.845 -19.555 ;
        RECT 237.155 -19.885 237.485 -19.555 ;
        RECT 235.795 -19.885 236.125 -19.555 ;
        RECT 234.435 -19.885 234.765 -19.555 ;
        RECT 233.075 -19.885 233.405 -19.555 ;
        RECT 231.715 -19.885 232.045 -19.555 ;
        RECT 227.635 -19.885 227.965 -19.555 ;
        RECT 224.915 -19.885 225.245 -19.555 ;
        RECT 223.555 -19.885 223.885 -19.555 ;
        RECT 222.195 -19.885 222.525 -19.555 ;
        RECT 220.835 -19.885 221.165 -19.555 ;
        RECT 219.475 -19.885 219.805 -19.555 ;
        RECT 218.115 -19.885 218.445 -19.555 ;
        RECT 216.755 -19.885 217.085 -19.555 ;
        RECT 212.675 -19.885 213.005 -19.555 ;
        RECT 209.955 -19.885 210.285 -19.555 ;
        RECT 208.595 -19.885 208.925 -19.555 ;
        RECT 207.235 -19.885 207.565 -19.555 ;
        RECT 205.875 -19.885 206.205 -19.555 ;
        RECT 204.515 -19.885 204.845 -19.555 ;
        RECT 203.155 -19.885 203.485 -19.555 ;
        RECT 201.795 -19.885 202.125 -19.555 ;
        RECT 197.715 -19.885 198.045 -19.555 ;
        RECT 194.995 -19.885 195.325 -19.555 ;
        RECT 193.635 -19.885 193.965 -19.555 ;
        RECT 192.275 -19.885 192.605 -19.555 ;
        RECT 190.915 -19.885 191.245 -19.555 ;
        RECT 189.555 -19.885 189.885 -19.555 ;
        RECT 188.195 -19.885 188.525 -19.555 ;
        RECT 186.835 -19.885 187.165 -19.555 ;
        RECT 182.755 -19.885 183.085 -19.555 ;
        RECT 180.035 -19.885 180.365 -19.555 ;
        RECT 178.675 -19.885 179.005 -19.555 ;
        RECT 177.315 -19.885 177.645 -19.555 ;
        RECT 175.955 -19.885 176.285 -19.555 ;
        RECT 174.595 -19.885 174.925 -19.555 ;
        RECT 173.235 -19.885 173.565 -19.555 ;
        RECT 171.875 -19.885 172.205 -19.555 ;
        RECT 167.795 -19.885 168.125 -19.555 ;
        RECT 165.075 -19.885 165.405 -19.555 ;
        RECT 163.715 -19.885 164.045 -19.555 ;
        RECT 162.355 -19.885 162.685 -19.555 ;
        RECT 160.995 -19.885 161.325 -19.555 ;
        RECT 159.635 -19.885 159.965 -19.555 ;
        RECT 158.275 -19.885 158.605 -19.555 ;
        RECT 156.915 -19.885 157.245 -19.555 ;
        RECT 152.835 -19.885 153.165 -19.555 ;
        RECT 150.115 -19.885 150.445 -19.555 ;
        RECT 148.755 -19.885 149.085 -19.555 ;
        RECT 147.395 -19.885 147.725 -19.555 ;
        RECT 146.035 -19.885 146.365 -19.555 ;
        RECT 144.675 -19.885 145.005 -19.555 ;
        RECT 143.315 -19.885 143.645 -19.555 ;
        RECT 141.955 -19.885 142.285 -19.555 ;
        RECT 136.515 -19.885 136.845 -19.555 ;
        RECT 135.155 -19.885 135.485 -19.555 ;
        RECT 133.795 -19.885 134.125 -19.555 ;
        RECT 132.435 -19.885 132.765 -19.555 ;
        RECT 131.075 -19.885 131.405 -19.555 ;
        RECT 129.715 -19.885 130.045 -19.555 ;
        RECT 128.355 -19.885 128.685 -19.555 ;
        RECT 126.995 -19.885 127.325 -19.555 ;
        RECT 121.555 -19.885 121.885 -19.555 ;
        RECT 120.195 -19.885 120.525 -19.555 ;
        RECT 118.835 -19.885 119.165 -19.555 ;
        RECT 117.475 -19.885 117.805 -19.555 ;
        RECT 116.115 -19.885 116.445 -19.555 ;
        RECT 114.755 -19.885 115.085 -19.555 ;
        RECT 113.395 -19.885 113.725 -19.555 ;
        RECT 112.035 -19.885 112.365 -19.555 ;
        RECT 106.595 -19.885 106.925 -19.555 ;
        RECT 105.235 -19.885 105.565 -19.555 ;
        RECT 103.875 -19.885 104.205 -19.555 ;
        RECT 102.515 -19.885 102.845 -19.555 ;
        RECT 101.155 -19.885 101.485 -19.555 ;
        RECT 99.795 -19.885 100.125 -19.555 ;
        RECT 98.435 -19.885 98.765 -19.555 ;
        RECT 97.075 -19.885 97.405 -19.555 ;
        RECT 91.635 -19.885 91.965 -19.555 ;
        RECT 90.275 -19.885 90.605 -19.555 ;
        RECT 88.915 -19.885 89.245 -19.555 ;
        RECT 87.555 -19.885 87.885 -19.555 ;
        RECT 86.195 -19.885 86.525 -19.555 ;
        RECT 84.835 -19.885 85.165 -19.555 ;
        RECT 83.475 -19.885 83.805 -19.555 ;
        RECT 82.115 -19.885 82.445 -19.555 ;
        RECT 76.675 -19.885 77.005 -19.555 ;
        RECT 75.315 -19.885 75.645 -19.555 ;
        RECT 73.955 -19.885 74.285 -19.555 ;
        RECT 72.595 -19.885 72.925 -19.555 ;
        RECT 71.235 -19.885 71.565 -19.555 ;
        RECT 69.875 -19.885 70.205 -19.555 ;
        RECT 68.515 -19.885 68.845 -19.555 ;
        RECT 67.155 -19.885 67.485 -19.555 ;
        RECT 61.715 -19.885 62.045 -19.555 ;
        RECT 60.355 -19.885 60.685 -19.555 ;
        RECT 58.995 -19.885 59.325 -19.555 ;
        RECT 57.635 -19.885 57.965 -19.555 ;
        RECT 56.275 -19.885 56.605 -19.555 ;
        RECT 54.915 -19.885 55.245 -19.555 ;
        RECT 53.555 -19.885 53.885 -19.555 ;
        RECT 52.195 -19.885 52.525 -19.555 ;
        RECT 46.755 -19.885 47.085 -19.555 ;
        RECT 45.395 -19.885 45.725 -19.555 ;
        RECT 44.035 -19.885 44.365 -19.555 ;
        RECT 42.675 -19.885 43.005 -19.555 ;
        RECT 41.315 -19.885 41.645 -19.555 ;
        RECT 39.955 -19.885 40.285 -19.555 ;
        RECT 38.595 -19.885 38.925 -19.555 ;
        RECT 37.235 -19.885 37.565 -19.555 ;
        RECT 31.795 -19.885 32.125 -19.555 ;
        RECT 30.435 -19.885 30.765 -19.555 ;
        RECT 29.075 -19.885 29.405 -19.555 ;
        RECT 27.715 -19.885 28.045 -19.555 ;
        RECT 26.355 -19.885 26.685 -19.555 ;
        RECT 24.995 -19.885 25.325 -19.555 ;
        RECT 23.635 -19.885 23.965 -19.555 ;
        RECT 22.275 -19.885 22.605 -19.555 ;
        RECT 16.835 -19.885 17.165 -19.555 ;
        RECT 15.475 -19.885 15.805 -19.555 ;
        RECT 14.115 -19.885 14.445 -19.555 ;
        RECT 12.755 -19.885 13.085 -19.555 ;
        RECT 11.395 -19.885 11.725 -19.555 ;
        RECT 10.035 -19.885 10.365 -19.555 ;
        RECT 8.675 -19.885 9.005 -19.555 ;
        RECT 7.315 -19.885 7.645 -19.555 ;
        RECT 3.235 -19.885 3.565 -19.555 ;
        RECT 1.875 -19.885 2.205 -19.555 ;
        RECT 0.515 -19.885 0.845 -19.555 ;
        RECT -0.845 -19.885 -0.515 -19.555 ;
        RECT 924.285 -19.88 954.88 -19.56 ;
        RECT 953.875 -19.885 954.205 -19.555 ;
        RECT 952.515 -19.885 952.845 -19.555 ;
        RECT 951.155 -19.885 951.485 -19.555 ;
        RECT 949.795 -19.885 950.125 -19.555 ;
        RECT 948.435 -19.885 948.765 -19.555 ;
        RECT 947.075 -19.885 947.405 -19.555 ;
        RECT 945.715 -19.885 946.045 -19.555 ;
        RECT 942.995 -19.885 943.325 -19.555 ;
        RECT 940.275 -19.885 940.605 -19.555 ;
        RECT 938.915 -19.885 939.245 -19.555 ;
        RECT 937.555 -19.885 937.885 -19.555 ;
        RECT 936.195 -19.885 936.525 -19.555 ;
        RECT 934.835 -19.885 935.165 -19.555 ;
        RECT 933.475 -19.885 933.805 -19.555 ;
        RECT 932.115 -19.885 932.445 -19.555 ;
        RECT 930.755 -19.885 931.085 -19.555 ;
        RECT 928.035 -19.885 928.365 -19.555 ;
        RECT 925.315 -19.885 925.645 -19.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 919.88 -29.4 926.32 -29.08 ;
        RECT 925.315 -29.405 925.645 -29.075 ;
        RECT 923.955 -29.405 924.285 -29.075 ;
        RECT 922.595 -29.405 922.925 -29.075 ;
        RECT 921.235 -29.405 921.565 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 915.8 -23.96 927 -23.64 ;
        RECT 925.315 -23.965 925.645 -23.635 ;
        RECT 923.955 -23.965 924.285 -23.635 ;
        RECT 922.595 -23.965 922.925 -23.635 ;
        RECT 921.235 -23.965 921.565 -23.635 ;
        RECT 919.875 -23.965 920.205 -23.635 ;
        RECT 917.155 -23.965 917.485 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 916.48 -28.04 927 -27.72 ;
        RECT 925.315 -28.045 925.645 -27.715 ;
        RECT 923.955 -28.045 924.285 -27.715 ;
        RECT 922.595 -28.045 922.925 -27.715 ;
        RECT 921.235 -28.045 921.565 -27.715 ;
        RECT 917.155 -28.045 917.485 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 926.675 -34.845 927.005 -34.515 ;
        RECT 919.88 -34.84 927.005 -34.52 ;
        RECT 925.315 -34.845 925.645 -34.515 ;
        RECT 923.955 -34.845 924.285 -34.515 ;
        RECT 922.595 -34.845 922.925 -34.515 ;
        RECT 921.235 -34.845 921.565 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 919.88 -26.68 930.4 -26.36 ;
        RECT 928.035 -26.685 928.365 -26.355 ;
        RECT 925.315 -26.685 925.645 -26.355 ;
        RECT 923.955 -26.685 924.285 -26.355 ;
        RECT 922.595 -26.685 922.925 -26.355 ;
        RECT 921.235 -26.685 921.565 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 930.755 -23.96 941.28 -23.64 ;
        RECT 940.275 -23.965 940.605 -23.635 ;
        RECT 938.915 -23.965 939.245 -23.635 ;
        RECT 937.555 -23.965 937.885 -23.635 ;
        RECT 936.195 -23.965 936.525 -23.635 ;
        RECT 934.835 -23.965 935.165 -23.635 ;
        RECT 932.115 -23.965 932.445 -23.635 ;
        RECT 930.755 -23.965 931.085 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 934.84 -34.84 944 -34.52 ;
        RECT 942.995 -34.845 943.325 -34.515 ;
        RECT 941.635 -34.845 941.965 -34.515 ;
        RECT 940.275 -34.845 940.605 -34.515 ;
        RECT 938.915 -34.845 939.245 -34.515 ;
        RECT 937.555 -34.845 937.885 -34.515 ;
        RECT 936.195 -34.845 936.525 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.875 -29.4 687.64 -29.08 ;
        RECT 685.955 -29.405 686.285 -29.075 ;
        RECT 684.595 -29.405 684.925 -29.075 ;
        RECT 683.235 -29.405 683.565 -29.075 ;
        RECT 681.875 -29.405 682.205 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.12 -23.96 688.32 -23.64 ;
        RECT 685.955 -23.965 686.285 -23.635 ;
        RECT 684.595 -23.965 684.925 -23.635 ;
        RECT 683.235 -23.965 683.565 -23.635 ;
        RECT 681.875 -23.965 682.205 -23.635 ;
        RECT 679.155 -23.965 679.485 -23.635 ;
        RECT 677.795 -23.965 678.125 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.8 -28.04 688.32 -27.72 ;
        RECT 685.955 -28.045 686.285 -27.715 ;
        RECT 684.595 -28.045 684.925 -27.715 ;
        RECT 683.235 -28.045 683.565 -27.715 ;
        RECT 681.875 -28.045 682.205 -27.715 ;
        RECT 679.155 -28.045 679.485 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.875 -34.84 688.32 -34.52 ;
        RECT 687.315 -34.845 687.645 -34.515 ;
        RECT 685.955 -34.845 686.285 -34.515 ;
        RECT 684.595 -34.845 684.925 -34.515 ;
        RECT 683.235 -34.845 683.565 -34.515 ;
        RECT 681.875 -34.845 682.205 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.875 -26.68 692.4 -26.36 ;
        RECT 690.035 -26.685 690.365 -26.355 ;
        RECT 685.955 -26.685 686.285 -26.355 ;
        RECT 684.595 -26.685 684.925 -26.355 ;
        RECT 683.235 -26.685 683.565 -26.355 ;
        RECT 681.875 -26.685 682.205 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.16 -29.4 702.6 -29.08 ;
        RECT 700.915 -29.405 701.245 -29.075 ;
        RECT 699.555 -29.405 699.885 -29.075 ;
        RECT 698.195 -29.405 698.525 -29.075 ;
        RECT 696.835 -29.405 697.165 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.08 -23.96 703.28 -23.64 ;
        RECT 700.915 -23.965 701.245 -23.635 ;
        RECT 699.555 -23.965 699.885 -23.635 ;
        RECT 698.195 -23.965 698.525 -23.635 ;
        RECT 696.835 -23.965 697.165 -23.635 ;
        RECT 692.755 -23.965 693.085 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.76 -28.04 703.28 -27.72 ;
        RECT 700.915 -28.045 701.245 -27.715 ;
        RECT 699.555 -28.045 699.885 -27.715 ;
        RECT 698.195 -28.045 698.525 -27.715 ;
        RECT 696.835 -28.045 697.165 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.16 -34.84 703.28 -34.52 ;
        RECT 702.275 -34.845 702.605 -34.515 ;
        RECT 700.915 -34.845 701.245 -34.515 ;
        RECT 699.555 -34.845 699.885 -34.515 ;
        RECT 698.195 -34.845 698.525 -34.515 ;
        RECT 696.835 -34.845 697.165 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.16 -26.68 707.36 -26.36 ;
        RECT 704.995 -26.685 705.325 -26.355 ;
        RECT 700.915 -26.685 701.245 -26.355 ;
        RECT 699.555 -26.685 699.885 -26.355 ;
        RECT 698.195 -26.685 698.525 -26.355 ;
        RECT 696.835 -26.685 697.165 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.12 -29.4 717.56 -29.08 ;
        RECT 715.875 -29.405 716.205 -29.075 ;
        RECT 714.515 -29.405 714.845 -29.075 ;
        RECT 713.155 -29.405 713.485 -29.075 ;
        RECT 711.795 -29.405 712.125 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.04 -23.96 718.24 -23.64 ;
        RECT 715.875 -23.965 716.205 -23.635 ;
        RECT 714.515 -23.965 714.845 -23.635 ;
        RECT 713.155 -23.965 713.485 -23.635 ;
        RECT 711.795 -23.965 712.125 -23.635 ;
        RECT 707.715 -23.965 708.045 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.72 -28.04 718.24 -27.72 ;
        RECT 715.875 -28.045 716.205 -27.715 ;
        RECT 714.515 -28.045 714.845 -27.715 ;
        RECT 713.155 -28.045 713.485 -27.715 ;
        RECT 711.795 -28.045 712.125 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.12 -34.84 718.24 -34.52 ;
        RECT 717.235 -34.845 717.565 -34.515 ;
        RECT 715.875 -34.845 716.205 -34.515 ;
        RECT 714.515 -34.845 714.845 -34.515 ;
        RECT 713.155 -34.845 713.485 -34.515 ;
        RECT 711.795 -34.845 712.125 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.12 -26.68 722.32 -26.36 ;
        RECT 719.955 -26.685 720.285 -26.355 ;
        RECT 715.875 -26.685 716.205 -26.355 ;
        RECT 714.515 -26.685 714.845 -26.355 ;
        RECT 713.155 -26.685 713.485 -26.355 ;
        RECT 711.795 -26.685 712.125 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.08 -29.4 732.52 -29.08 ;
        RECT 730.835 -29.405 731.165 -29.075 ;
        RECT 729.475 -29.405 729.805 -29.075 ;
        RECT 728.115 -29.405 728.445 -29.075 ;
        RECT 726.755 -29.405 727.085 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 722 -23.96 733.2 -23.64 ;
        RECT 730.835 -23.965 731.165 -23.635 ;
        RECT 729.475 -23.965 729.805 -23.635 ;
        RECT 728.115 -23.965 728.445 -23.635 ;
        RECT 726.755 -23.965 727.085 -23.635 ;
        RECT 722.675 -23.965 723.005 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 722.68 -28.04 733.2 -27.72 ;
        RECT 730.835 -28.045 731.165 -27.715 ;
        RECT 729.475 -28.045 729.805 -27.715 ;
        RECT 728.115 -28.045 728.445 -27.715 ;
        RECT 726.755 -28.045 727.085 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.08 -34.84 733.2 -34.52 ;
        RECT 732.195 -34.845 732.525 -34.515 ;
        RECT 730.835 -34.845 731.165 -34.515 ;
        RECT 729.475 -34.845 729.805 -34.515 ;
        RECT 728.115 -34.845 728.445 -34.515 ;
        RECT 726.755 -34.845 727.085 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.08 -26.68 736.6 -26.36 ;
        RECT 734.915 -26.685 735.245 -26.355 ;
        RECT 730.835 -26.685 731.165 -26.355 ;
        RECT 729.475 -26.685 729.805 -26.355 ;
        RECT 728.115 -26.685 728.445 -26.355 ;
        RECT 726.755 -26.685 727.085 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.04 -29.4 747.48 -29.08 ;
        RECT 745.795 -29.405 746.125 -29.075 ;
        RECT 744.435 -29.405 744.765 -29.075 ;
        RECT 743.075 -29.405 743.405 -29.075 ;
        RECT 741.715 -29.405 742.045 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.96 -23.96 748.16 -23.64 ;
        RECT 745.795 -23.965 746.125 -23.635 ;
        RECT 744.435 -23.965 744.765 -23.635 ;
        RECT 743.075 -23.965 743.405 -23.635 ;
        RECT 741.715 -23.965 742.045 -23.635 ;
        RECT 737.635 -23.965 737.965 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 737.64 -28.04 748.16 -27.72 ;
        RECT 745.795 -28.045 746.125 -27.715 ;
        RECT 744.435 -28.045 744.765 -27.715 ;
        RECT 743.075 -28.045 743.405 -27.715 ;
        RECT 741.715 -28.045 742.045 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.04 -34.84 748.16 -34.52 ;
        RECT 747.155 -34.845 747.485 -34.515 ;
        RECT 745.795 -34.845 746.125 -34.515 ;
        RECT 744.435 -34.845 744.765 -34.515 ;
        RECT 743.075 -34.845 743.405 -34.515 ;
        RECT 741.715 -34.845 742.045 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.04 -26.68 751.56 -26.36 ;
        RECT 749.875 -26.685 750.205 -26.355 ;
        RECT 745.795 -26.685 746.125 -26.355 ;
        RECT 744.435 -26.685 744.765 -26.355 ;
        RECT 743.075 -26.685 743.405 -26.355 ;
        RECT 741.715 -26.685 742.045 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 756 -29.4 762.44 -29.08 ;
        RECT 760.755 -29.405 761.085 -29.075 ;
        RECT 759.395 -29.405 759.725 -29.075 ;
        RECT 758.035 -29.405 758.365 -29.075 ;
        RECT 756.675 -29.405 757.005 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.92 -23.96 763.12 -23.64 ;
        RECT 760.755 -23.965 761.085 -23.635 ;
        RECT 759.395 -23.965 759.725 -23.635 ;
        RECT 758.035 -23.965 758.365 -23.635 ;
        RECT 756.675 -23.965 757.005 -23.635 ;
        RECT 752.595 -23.965 752.925 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 752.6 -28.04 763.12 -27.72 ;
        RECT 760.755 -28.045 761.085 -27.715 ;
        RECT 759.395 -28.045 759.725 -27.715 ;
        RECT 758.035 -28.045 758.365 -27.715 ;
        RECT 756.675 -28.045 757.005 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 756 -34.84 763.12 -34.52 ;
        RECT 762.115 -34.845 762.445 -34.515 ;
        RECT 760.755 -34.845 761.085 -34.515 ;
        RECT 759.395 -34.845 759.725 -34.515 ;
        RECT 758.035 -34.845 758.365 -34.515 ;
        RECT 756.675 -34.845 757.005 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 756 -26.68 766.52 -26.36 ;
        RECT 764.835 -26.685 765.165 -26.355 ;
        RECT 760.755 -26.685 761.085 -26.355 ;
        RECT 759.395 -26.685 759.725 -26.355 ;
        RECT 758.035 -26.685 758.365 -26.355 ;
        RECT 756.675 -26.685 757.005 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 770.96 -29.4 777.4 -29.08 ;
        RECT 775.715 -29.405 776.045 -29.075 ;
        RECT 774.355 -29.405 774.685 -29.075 ;
        RECT 772.995 -29.405 773.325 -29.075 ;
        RECT 771.635 -29.405 771.965 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.955 -18.525 652.285 -18.195 ;
        RECT 650.595 -18.525 650.925 -18.195 ;
        RECT 649.235 -18.525 649.565 -18.195 ;
        RECT 647.875 -18.525 648.205 -18.195 ;
        RECT 645.155 -18.525 645.485 -18.195 ;
        RECT 643.795 -18.525 644.125 -18.195 ;
        RECT 642.435 -18.525 642.765 -18.195 ;
        RECT 641.075 -18.525 641.405 -18.195 ;
        RECT 639.715 -18.525 640.045 -18.195 ;
        RECT 638.355 -18.525 638.685 -18.195 ;
        RECT 636.995 -18.525 637.325 -18.195 ;
        RECT 635.635 -18.525 635.965 -18.195 ;
        RECT 634.275 -18.525 634.605 -18.195 ;
        RECT 632.915 -18.525 633.245 -18.195 ;
        RECT 630.195 -18.525 630.525 -18.195 ;
        RECT 628.835 -18.525 629.165 -18.195 ;
        RECT 627.475 -18.525 627.805 -18.195 ;
        RECT 626.115 -18.525 626.445 -18.195 ;
        RECT 624.755 -18.525 625.085 -18.195 ;
        RECT 623.395 -18.525 623.725 -18.195 ;
        RECT 622.035 -18.525 622.365 -18.195 ;
        RECT 620.675 -18.525 621.005 -18.195 ;
        RECT 619.315 -18.525 619.645 -18.195 ;
        RECT 617.955 -18.525 618.285 -18.195 ;
        RECT 615.235 -18.525 615.565 -18.195 ;
        RECT 613.875 -18.525 614.205 -18.195 ;
        RECT 612.515 -18.525 612.845 -18.195 ;
        RECT 611.155 -18.525 611.485 -18.195 ;
        RECT 609.795 -18.525 610.125 -18.195 ;
        RECT 608.435 -18.525 608.765 -18.195 ;
        RECT 607.075 -18.525 607.405 -18.195 ;
        RECT 605.715 -18.525 606.045 -18.195 ;
        RECT 604.355 -18.525 604.685 -18.195 ;
        RECT 602.995 -18.525 603.325 -18.195 ;
        RECT 600.275 -18.525 600.605 -18.195 ;
        RECT 598.915 -18.525 599.245 -18.195 ;
        RECT 597.555 -18.525 597.885 -18.195 ;
        RECT 596.195 -18.525 596.525 -18.195 ;
        RECT 594.835 -18.525 595.165 -18.195 ;
        RECT 593.475 -18.525 593.805 -18.195 ;
        RECT 592.115 -18.525 592.445 -18.195 ;
        RECT 590.755 -18.525 591.085 -18.195 ;
        RECT 589.395 -18.525 589.725 -18.195 ;
        RECT 588.035 -18.525 588.365 -18.195 ;
        RECT 585.315 -18.525 585.645 -18.195 ;
        RECT 583.955 -18.525 584.285 -18.195 ;
        RECT 582.595 -18.525 582.925 -18.195 ;
        RECT 581.235 -18.525 581.565 -18.195 ;
        RECT 579.875 -18.525 580.205 -18.195 ;
        RECT 578.515 -18.525 578.845 -18.195 ;
        RECT 577.155 -18.525 577.485 -18.195 ;
        RECT 575.795 -18.525 576.125 -18.195 ;
        RECT 574.435 -18.525 574.765 -18.195 ;
        RECT 570.355 -18.525 570.685 -18.195 ;
        RECT 568.995 -18.525 569.325 -18.195 ;
        RECT 567.635 -18.525 567.965 -18.195 ;
        RECT 566.275 -18.525 566.605 -18.195 ;
        RECT 564.915 -18.525 565.245 -18.195 ;
        RECT 563.555 -18.525 563.885 -18.195 ;
        RECT 562.195 -18.525 562.525 -18.195 ;
        RECT 560.835 -18.525 561.165 -18.195 ;
        RECT 559.475 -18.525 559.805 -18.195 ;
        RECT 555.395 -18.525 555.725 -18.195 ;
        RECT 554.035 -18.525 554.365 -18.195 ;
        RECT 552.675 -18.525 553.005 -18.195 ;
        RECT 551.315 -18.525 551.645 -18.195 ;
        RECT 549.955 -18.525 550.285 -18.195 ;
        RECT 548.595 -18.525 548.925 -18.195 ;
        RECT 547.235 -18.525 547.565 -18.195 ;
        RECT 545.875 -18.525 546.205 -18.195 ;
        RECT 544.515 -18.525 544.845 -18.195 ;
        RECT 540.435 -18.525 540.765 -18.195 ;
        RECT 539.075 -18.525 539.405 -18.195 ;
        RECT 537.715 -18.525 538.045 -18.195 ;
        RECT 536.355 -18.525 536.685 -18.195 ;
        RECT 534.995 -18.525 535.325 -18.195 ;
        RECT 533.635 -18.525 533.965 -18.195 ;
        RECT 532.275 -18.525 532.605 -18.195 ;
        RECT 530.915 -18.525 531.245 -18.195 ;
        RECT 529.555 -18.525 529.885 -18.195 ;
        RECT 525.475 -18.525 525.805 -18.195 ;
        RECT 524.115 -18.525 524.445 -18.195 ;
        RECT 522.755 -18.525 523.085 -18.195 ;
        RECT 521.395 -18.525 521.725 -18.195 ;
        RECT 520.035 -18.525 520.365 -18.195 ;
        RECT 518.675 -18.525 519.005 -18.195 ;
        RECT 517.315 -18.525 517.645 -18.195 ;
        RECT 515.955 -18.525 516.285 -18.195 ;
        RECT 514.595 -18.525 514.925 -18.195 ;
        RECT 510.515 -18.525 510.845 -18.195 ;
        RECT 509.155 -18.525 509.485 -18.195 ;
        RECT 507.795 -18.525 508.125 -18.195 ;
        RECT 506.435 -18.525 506.765 -18.195 ;
        RECT 505.075 -18.525 505.405 -18.195 ;
        RECT 503.715 -18.525 504.045 -18.195 ;
        RECT 502.355 -18.525 502.685 -18.195 ;
        RECT 500.995 -18.525 501.325 -18.195 ;
        RECT 499.635 -18.525 499.965 -18.195 ;
        RECT 495.555 -18.525 495.885 -18.195 ;
        RECT 494.195 -18.525 494.525 -18.195 ;
        RECT 492.835 -18.525 493.165 -18.195 ;
        RECT 491.475 -18.525 491.805 -18.195 ;
        RECT 490.115 -18.525 490.445 -18.195 ;
        RECT 488.755 -18.525 489.085 -18.195 ;
        RECT 487.395 -18.525 487.725 -18.195 ;
        RECT 486.035 -18.525 486.365 -18.195 ;
        RECT 484.675 -18.525 485.005 -18.195 ;
        RECT 480.595 -18.525 480.925 -18.195 ;
        RECT 479.235 -18.525 479.565 -18.195 ;
        RECT 477.875 -18.525 478.205 -18.195 ;
        RECT 476.515 -18.525 476.845 -18.195 ;
        RECT 475.155 -18.525 475.485 -18.195 ;
        RECT 473.795 -18.525 474.125 -18.195 ;
        RECT 472.435 -18.525 472.765 -18.195 ;
        RECT 471.075 -18.525 471.405 -18.195 ;
        RECT 469.715 -18.525 470.045 -18.195 ;
        RECT 465.635 -18.525 465.965 -18.195 ;
        RECT 464.275 -18.525 464.605 -18.195 ;
        RECT 462.915 -18.525 463.245 -18.195 ;
        RECT 461.555 -18.525 461.885 -18.195 ;
        RECT 460.195 -18.525 460.525 -18.195 ;
        RECT 458.835 -18.525 459.165 -18.195 ;
        RECT 457.475 -18.525 457.805 -18.195 ;
        RECT 456.115 -18.525 456.445 -18.195 ;
        RECT 454.755 -18.525 455.085 -18.195 ;
        RECT 450.675 -18.525 451.005 -18.195 ;
        RECT 449.315 -18.525 449.645 -18.195 ;
        RECT 447.955 -18.525 448.285 -18.195 ;
        RECT 446.595 -18.525 446.925 -18.195 ;
        RECT 445.235 -18.525 445.565 -18.195 ;
        RECT 443.875 -18.525 444.205 -18.195 ;
        RECT 442.515 -18.525 442.845 -18.195 ;
        RECT 441.155 -18.525 441.485 -18.195 ;
        RECT 439.795 -18.525 440.125 -18.195 ;
        RECT 435.715 -18.525 436.045 -18.195 ;
        RECT 434.355 -18.525 434.685 -18.195 ;
        RECT 432.995 -18.525 433.325 -18.195 ;
        RECT 431.635 -18.525 431.965 -18.195 ;
        RECT 430.275 -18.525 430.605 -18.195 ;
        RECT 428.915 -18.525 429.245 -18.195 ;
        RECT 427.555 -18.525 427.885 -18.195 ;
        RECT 426.195 -18.525 426.525 -18.195 ;
        RECT 424.835 -18.525 425.165 -18.195 ;
        RECT 422.115 -18.525 422.445 -18.195 ;
        RECT 420.755 -18.525 421.085 -18.195 ;
        RECT 419.395 -18.525 419.725 -18.195 ;
        RECT 418.035 -18.525 418.365 -18.195 ;
        RECT 416.675 -18.525 417.005 -18.195 ;
        RECT 415.315 -18.525 415.645 -18.195 ;
        RECT 413.955 -18.525 414.285 -18.195 ;
        RECT 412.595 -18.525 412.925 -18.195 ;
        RECT 411.235 -18.525 411.565 -18.195 ;
        RECT 409.875 -18.525 410.205 -18.195 ;
        RECT 407.155 -18.525 407.485 -18.195 ;
        RECT 405.795 -18.525 406.125 -18.195 ;
        RECT 404.435 -18.525 404.765 -18.195 ;
        RECT 403.075 -18.525 403.405 -18.195 ;
        RECT 401.715 -18.525 402.045 -18.195 ;
        RECT 400.355 -18.525 400.685 -18.195 ;
        RECT 398.995 -18.525 399.325 -18.195 ;
        RECT 397.635 -18.525 397.965 -18.195 ;
        RECT 396.275 -18.525 396.605 -18.195 ;
        RECT 394.915 -18.525 395.245 -18.195 ;
        RECT 392.195 -18.525 392.525 -18.195 ;
        RECT 390.835 -18.525 391.165 -18.195 ;
        RECT 389.475 -18.525 389.805 -18.195 ;
        RECT 388.115 -18.525 388.445 -18.195 ;
        RECT 386.755 -18.525 387.085 -18.195 ;
        RECT 385.395 -18.525 385.725 -18.195 ;
        RECT 384.035 -18.525 384.365 -18.195 ;
        RECT 382.675 -18.525 383.005 -18.195 ;
        RECT 381.315 -18.525 381.645 -18.195 ;
        RECT 379.955 -18.525 380.285 -18.195 ;
        RECT 377.235 -18.525 377.565 -18.195 ;
        RECT 375.875 -18.525 376.205 -18.195 ;
        RECT 374.515 -18.525 374.845 -18.195 ;
        RECT 373.155 -18.525 373.485 -18.195 ;
        RECT 371.795 -18.525 372.125 -18.195 ;
        RECT 370.435 -18.525 370.765 -18.195 ;
        RECT 369.075 -18.525 369.405 -18.195 ;
        RECT 367.715 -18.525 368.045 -18.195 ;
        RECT 366.355 -18.525 366.685 -18.195 ;
        RECT 364.995 -18.525 365.325 -18.195 ;
        RECT 362.275 -18.525 362.605 -18.195 ;
        RECT 360.915 -18.525 361.245 -18.195 ;
        RECT 359.555 -18.525 359.885 -18.195 ;
        RECT 358.195 -18.525 358.525 -18.195 ;
        RECT 356.835 -18.525 357.165 -18.195 ;
        RECT 355.475 -18.525 355.805 -18.195 ;
        RECT 354.115 -18.525 354.445 -18.195 ;
        RECT 352.755 -18.525 353.085 -18.195 ;
        RECT 351.395 -18.525 351.725 -18.195 ;
        RECT 350.035 -18.525 350.365 -18.195 ;
        RECT 347.315 -18.525 347.645 -18.195 ;
        RECT 345.955 -18.525 346.285 -18.195 ;
        RECT 344.595 -18.525 344.925 -18.195 ;
        RECT 343.235 -18.525 343.565 -18.195 ;
        RECT 341.875 -18.525 342.205 -18.195 ;
        RECT 340.515 -18.525 340.845 -18.195 ;
        RECT 339.155 -18.525 339.485 -18.195 ;
        RECT 337.795 -18.525 338.125 -18.195 ;
        RECT 336.435 -18.525 336.765 -18.195 ;
        RECT 335.075 -18.525 335.405 -18.195 ;
        RECT 332.355 -18.525 332.685 -18.195 ;
        RECT 330.995 -18.525 331.325 -18.195 ;
        RECT 329.635 -18.525 329.965 -18.195 ;
        RECT 328.275 -18.525 328.605 -18.195 ;
        RECT 326.915 -18.525 327.245 -18.195 ;
        RECT 325.555 -18.525 325.885 -18.195 ;
        RECT 324.195 -18.525 324.525 -18.195 ;
        RECT 322.835 -18.525 323.165 -18.195 ;
        RECT 321.475 -18.525 321.805 -18.195 ;
        RECT 320.115 -18.525 320.445 -18.195 ;
        RECT 317.395 -18.525 317.725 -18.195 ;
        RECT 316.035 -18.525 316.365 -18.195 ;
        RECT 314.675 -18.525 315.005 -18.195 ;
        RECT 313.315 -18.525 313.645 -18.195 ;
        RECT 311.955 -18.525 312.285 -18.195 ;
        RECT 310.595 -18.525 310.925 -18.195 ;
        RECT 309.235 -18.525 309.565 -18.195 ;
        RECT 307.875 -18.525 308.205 -18.195 ;
        RECT 306.515 -18.525 306.845 -18.195 ;
        RECT 305.155 -18.525 305.485 -18.195 ;
        RECT 302.435 -18.525 302.765 -18.195 ;
        RECT 301.075 -18.525 301.405 -18.195 ;
        RECT 299.715 -18.525 300.045 -18.195 ;
        RECT 298.355 -18.525 298.685 -18.195 ;
        RECT 296.995 -18.525 297.325 -18.195 ;
        RECT 295.635 -18.525 295.965 -18.195 ;
        RECT 294.275 -18.525 294.605 -18.195 ;
        RECT 292.915 -18.525 293.245 -18.195 ;
        RECT 291.555 -18.525 291.885 -18.195 ;
        RECT 290.195 -18.525 290.525 -18.195 ;
        RECT 287.475 -18.525 287.805 -18.195 ;
        RECT 286.115 -18.525 286.445 -18.195 ;
        RECT 284.755 -18.525 285.085 -18.195 ;
        RECT 283.395 -18.525 283.725 -18.195 ;
        RECT 282.035 -18.525 282.365 -18.195 ;
        RECT 280.675 -18.525 281.005 -18.195 ;
        RECT 279.315 -18.525 279.645 -18.195 ;
        RECT 277.955 -18.525 278.285 -18.195 ;
        RECT 276.595 -18.525 276.925 -18.195 ;
        RECT 275.235 -18.525 275.565 -18.195 ;
        RECT 272.515 -18.525 272.845 -18.195 ;
        RECT 271.155 -18.525 271.485 -18.195 ;
        RECT 269.795 -18.525 270.125 -18.195 ;
        RECT 268.435 -18.525 268.765 -18.195 ;
        RECT 267.075 -18.525 267.405 -18.195 ;
        RECT 265.715 -18.525 266.045 -18.195 ;
        RECT 264.355 -18.525 264.685 -18.195 ;
        RECT 262.995 -18.525 263.325 -18.195 ;
        RECT 261.635 -18.525 261.965 -18.195 ;
        RECT 260.275 -18.525 260.605 -18.195 ;
        RECT 257.555 -18.525 257.885 -18.195 ;
        RECT 256.195 -18.525 256.525 -18.195 ;
        RECT 254.835 -18.525 255.165 -18.195 ;
        RECT 253.475 -18.525 253.805 -18.195 ;
        RECT 252.115 -18.525 252.445 -18.195 ;
        RECT 250.755 -18.525 251.085 -18.195 ;
        RECT 249.395 -18.525 249.725 -18.195 ;
        RECT 248.035 -18.525 248.365 -18.195 ;
        RECT 246.675 -18.525 247.005 -18.195 ;
        RECT 242.595 -18.525 242.925 -18.195 ;
        RECT 241.235 -18.525 241.565 -18.195 ;
        RECT 239.875 -18.525 240.205 -18.195 ;
        RECT 238.515 -18.525 238.845 -18.195 ;
        RECT 237.155 -18.525 237.485 -18.195 ;
        RECT 235.795 -18.525 236.125 -18.195 ;
        RECT 234.435 -18.525 234.765 -18.195 ;
        RECT 233.075 -18.525 233.405 -18.195 ;
        RECT 231.715 -18.525 232.045 -18.195 ;
        RECT 227.635 -18.525 227.965 -18.195 ;
        RECT 226.275 -18.525 226.605 -18.195 ;
        RECT 224.915 -18.525 225.245 -18.195 ;
        RECT 223.555 -18.525 223.885 -18.195 ;
        RECT 222.195 -18.525 222.525 -18.195 ;
        RECT 220.835 -18.525 221.165 -18.195 ;
        RECT 219.475 -18.525 219.805 -18.195 ;
        RECT 218.115 -18.525 218.445 -18.195 ;
        RECT 216.755 -18.525 217.085 -18.195 ;
        RECT 212.675 -18.525 213.005 -18.195 ;
        RECT 211.315 -18.525 211.645 -18.195 ;
        RECT 209.955 -18.525 210.285 -18.195 ;
        RECT 208.595 -18.525 208.925 -18.195 ;
        RECT 207.235 -18.525 207.565 -18.195 ;
        RECT 205.875 -18.525 206.205 -18.195 ;
        RECT 204.515 -18.525 204.845 -18.195 ;
        RECT 203.155 -18.525 203.485 -18.195 ;
        RECT 201.795 -18.525 202.125 -18.195 ;
        RECT 197.715 -18.525 198.045 -18.195 ;
        RECT 196.355 -18.525 196.685 -18.195 ;
        RECT 194.995 -18.525 195.325 -18.195 ;
        RECT 193.635 -18.525 193.965 -18.195 ;
        RECT 192.275 -18.525 192.605 -18.195 ;
        RECT 190.915 -18.525 191.245 -18.195 ;
        RECT 189.555 -18.525 189.885 -18.195 ;
        RECT 188.195 -18.525 188.525 -18.195 ;
        RECT 186.835 -18.525 187.165 -18.195 ;
        RECT 182.755 -18.525 183.085 -18.195 ;
        RECT 181.395 -18.525 181.725 -18.195 ;
        RECT 180.035 -18.525 180.365 -18.195 ;
        RECT 178.675 -18.525 179.005 -18.195 ;
        RECT 177.315 -18.525 177.645 -18.195 ;
        RECT 175.955 -18.525 176.285 -18.195 ;
        RECT 174.595 -18.525 174.925 -18.195 ;
        RECT 173.235 -18.525 173.565 -18.195 ;
        RECT 171.875 -18.525 172.205 -18.195 ;
        RECT 167.795 -18.525 168.125 -18.195 ;
        RECT 166.435 -18.525 166.765 -18.195 ;
        RECT 165.075 -18.525 165.405 -18.195 ;
        RECT 163.715 -18.525 164.045 -18.195 ;
        RECT 162.355 -18.525 162.685 -18.195 ;
        RECT 160.995 -18.525 161.325 -18.195 ;
        RECT 159.635 -18.525 159.965 -18.195 ;
        RECT 158.275 -18.525 158.605 -18.195 ;
        RECT 156.915 -18.525 157.245 -18.195 ;
        RECT 152.835 -18.525 153.165 -18.195 ;
        RECT 151.475 -18.525 151.805 -18.195 ;
        RECT 150.115 -18.525 150.445 -18.195 ;
        RECT 148.755 -18.525 149.085 -18.195 ;
        RECT 147.395 -18.525 147.725 -18.195 ;
        RECT 146.035 -18.525 146.365 -18.195 ;
        RECT 144.675 -18.525 145.005 -18.195 ;
        RECT 143.315 -18.525 143.645 -18.195 ;
        RECT 141.955 -18.525 142.285 -18.195 ;
        RECT 137.875 -18.525 138.205 -18.195 ;
        RECT 136.515 -18.525 136.845 -18.195 ;
        RECT 135.155 -18.525 135.485 -18.195 ;
        RECT 133.795 -18.525 134.125 -18.195 ;
        RECT 132.435 -18.525 132.765 -18.195 ;
        RECT 131.075 -18.525 131.405 -18.195 ;
        RECT 129.715 -18.525 130.045 -18.195 ;
        RECT 128.355 -18.525 128.685 -18.195 ;
        RECT 126.995 -18.525 127.325 -18.195 ;
        RECT 122.915 -18.525 123.245 -18.195 ;
        RECT 121.555 -18.525 121.885 -18.195 ;
        RECT 120.195 -18.525 120.525 -18.195 ;
        RECT 118.835 -18.525 119.165 -18.195 ;
        RECT 117.475 -18.525 117.805 -18.195 ;
        RECT 116.115 -18.525 116.445 -18.195 ;
        RECT 114.755 -18.525 115.085 -18.195 ;
        RECT 113.395 -18.525 113.725 -18.195 ;
        RECT 112.035 -18.525 112.365 -18.195 ;
        RECT 107.955 -18.525 108.285 -18.195 ;
        RECT 106.595 -18.525 106.925 -18.195 ;
        RECT 105.235 -18.525 105.565 -18.195 ;
        RECT 103.875 -18.525 104.205 -18.195 ;
        RECT 102.515 -18.525 102.845 -18.195 ;
        RECT 101.155 -18.525 101.485 -18.195 ;
        RECT 99.795 -18.525 100.125 -18.195 ;
        RECT 98.435 -18.525 98.765 -18.195 ;
        RECT 97.075 -18.525 97.405 -18.195 ;
        RECT 92.995 -18.525 93.325 -18.195 ;
        RECT 91.635 -18.525 91.965 -18.195 ;
        RECT 90.275 -18.525 90.605 -18.195 ;
        RECT 88.915 -18.525 89.245 -18.195 ;
        RECT 87.555 -18.525 87.885 -18.195 ;
        RECT 86.195 -18.525 86.525 -18.195 ;
        RECT 84.835 -18.525 85.165 -18.195 ;
        RECT 83.475 -18.525 83.805 -18.195 ;
        RECT 82.115 -18.525 82.445 -18.195 ;
        RECT 79.395 -18.525 79.725 -18.195 ;
        RECT 78.035 -18.525 78.365 -18.195 ;
        RECT 76.675 -18.525 77.005 -18.195 ;
        RECT 75.315 -18.525 75.645 -18.195 ;
        RECT 73.955 -18.525 74.285 -18.195 ;
        RECT 72.595 -18.525 72.925 -18.195 ;
        RECT 71.235 -18.525 71.565 -18.195 ;
        RECT 69.875 -18.525 70.205 -18.195 ;
        RECT 68.515 -18.525 68.845 -18.195 ;
        RECT 67.155 -18.525 67.485 -18.195 ;
        RECT 64.435 -18.525 64.765 -18.195 ;
        RECT 63.075 -18.525 63.405 -18.195 ;
        RECT 61.715 -18.525 62.045 -18.195 ;
        RECT 60.355 -18.525 60.685 -18.195 ;
        RECT 58.995 -18.525 59.325 -18.195 ;
        RECT 57.635 -18.525 57.965 -18.195 ;
        RECT 56.275 -18.525 56.605 -18.195 ;
        RECT 54.915 -18.525 55.245 -18.195 ;
        RECT 53.555 -18.525 53.885 -18.195 ;
        RECT 52.195 -18.525 52.525 -18.195 ;
        RECT 49.475 -18.525 49.805 -18.195 ;
        RECT 48.115 -18.525 48.445 -18.195 ;
        RECT 46.755 -18.525 47.085 -18.195 ;
        RECT 45.395 -18.525 45.725 -18.195 ;
        RECT 44.035 -18.525 44.365 -18.195 ;
        RECT 42.675 -18.525 43.005 -18.195 ;
        RECT 41.315 -18.525 41.645 -18.195 ;
        RECT 39.955 -18.525 40.285 -18.195 ;
        RECT 38.595 -18.525 38.925 -18.195 ;
        RECT 37.235 -18.525 37.565 -18.195 ;
        RECT 34.515 -18.525 34.845 -18.195 ;
        RECT 33.155 -18.525 33.485 -18.195 ;
        RECT 31.795 -18.525 32.125 -18.195 ;
        RECT 30.435 -18.525 30.765 -18.195 ;
        RECT 29.075 -18.525 29.405 -18.195 ;
        RECT 27.715 -18.525 28.045 -18.195 ;
        RECT 26.355 -18.525 26.685 -18.195 ;
        RECT 24.995 -18.525 25.325 -18.195 ;
        RECT 23.635 -18.525 23.965 -18.195 ;
        RECT 22.275 -18.525 22.605 -18.195 ;
        RECT 19.555 -18.525 19.885 -18.195 ;
        RECT 18.195 -18.525 18.525 -18.195 ;
        RECT 16.835 -18.525 17.165 -18.195 ;
        RECT 15.475 -18.525 15.805 -18.195 ;
        RECT 14.115 -18.525 14.445 -18.195 ;
        RECT 12.755 -18.525 13.085 -18.195 ;
        RECT 11.395 -18.525 11.725 -18.195 ;
        RECT 10.035 -18.525 10.365 -18.195 ;
        RECT 8.675 -18.525 9.005 -18.195 ;
        RECT 7.315 -18.525 7.645 -18.195 ;
        RECT 4.595 -18.525 4.925 -18.195 ;
        RECT 3.235 -18.525 3.565 -18.195 ;
        RECT 1.875 -18.525 2.205 -18.195 ;
        RECT 0.515 -18.525 0.845 -18.195 ;
        RECT -0.845 -18.525 -0.515 -18.195 ;
        RECT 777.075 -18.525 777.405 -18.195 ;
        RECT -1.52 -18.52 777.405 -18.2 ;
        RECT 775.715 -18.525 776.045 -18.195 ;
        RECT 774.355 -18.525 774.685 -18.195 ;
        RECT 772.995 -18.525 773.325 -18.195 ;
        RECT 771.635 -18.525 771.965 -18.195 ;
        RECT 770.275 -18.525 770.605 -18.195 ;
        RECT 768.915 -18.525 769.245 -18.195 ;
        RECT 767.555 -18.525 767.885 -18.195 ;
        RECT 764.835 -18.525 765.165 -18.195 ;
        RECT 763.475 -18.525 763.805 -18.195 ;
        RECT 762.115 -18.525 762.445 -18.195 ;
        RECT 760.755 -18.525 761.085 -18.195 ;
        RECT 759.395 -18.525 759.725 -18.195 ;
        RECT 758.035 -18.525 758.365 -18.195 ;
        RECT 756.675 -18.525 757.005 -18.195 ;
        RECT 755.315 -18.525 755.645 -18.195 ;
        RECT 753.955 -18.525 754.285 -18.195 ;
        RECT 752.595 -18.525 752.925 -18.195 ;
        RECT 749.875 -18.525 750.205 -18.195 ;
        RECT 748.515 -18.525 748.845 -18.195 ;
        RECT 747.155 -18.525 747.485 -18.195 ;
        RECT 745.795 -18.525 746.125 -18.195 ;
        RECT 744.435 -18.525 744.765 -18.195 ;
        RECT 743.075 -18.525 743.405 -18.195 ;
        RECT 741.715 -18.525 742.045 -18.195 ;
        RECT 740.355 -18.525 740.685 -18.195 ;
        RECT 738.995 -18.525 739.325 -18.195 ;
        RECT 737.635 -18.525 737.965 -18.195 ;
        RECT 734.915 -18.525 735.245 -18.195 ;
        RECT 733.555 -18.525 733.885 -18.195 ;
        RECT 732.195 -18.525 732.525 -18.195 ;
        RECT 730.835 -18.525 731.165 -18.195 ;
        RECT 729.475 -18.525 729.805 -18.195 ;
        RECT 728.115 -18.525 728.445 -18.195 ;
        RECT 726.755 -18.525 727.085 -18.195 ;
        RECT 725.395 -18.525 725.725 -18.195 ;
        RECT 724.035 -18.525 724.365 -18.195 ;
        RECT 722.675 -18.525 723.005 -18.195 ;
        RECT 719.955 -18.525 720.285 -18.195 ;
        RECT 718.595 -18.525 718.925 -18.195 ;
        RECT 717.235 -18.525 717.565 -18.195 ;
        RECT 715.875 -18.525 716.205 -18.195 ;
        RECT 714.515 -18.525 714.845 -18.195 ;
        RECT 713.155 -18.525 713.485 -18.195 ;
        RECT 711.795 -18.525 712.125 -18.195 ;
        RECT 710.435 -18.525 710.765 -18.195 ;
        RECT 709.075 -18.525 709.405 -18.195 ;
        RECT 707.715 -18.525 708.045 -18.195 ;
        RECT 704.995 -18.525 705.325 -18.195 ;
        RECT 703.635 -18.525 703.965 -18.195 ;
        RECT 702.275 -18.525 702.605 -18.195 ;
        RECT 700.915 -18.525 701.245 -18.195 ;
        RECT 699.555 -18.525 699.885 -18.195 ;
        RECT 698.195 -18.525 698.525 -18.195 ;
        RECT 696.835 -18.525 697.165 -18.195 ;
        RECT 695.475 -18.525 695.805 -18.195 ;
        RECT 694.115 -18.525 694.445 -18.195 ;
        RECT 692.755 -18.525 693.085 -18.195 ;
        RECT 690.035 -18.525 690.365 -18.195 ;
        RECT 688.675 -18.525 689.005 -18.195 ;
        RECT 687.315 -18.525 687.645 -18.195 ;
        RECT 685.955 -18.525 686.285 -18.195 ;
        RECT 684.595 -18.525 684.925 -18.195 ;
        RECT 683.235 -18.525 683.565 -18.195 ;
        RECT 681.875 -18.525 682.205 -18.195 ;
        RECT 680.515 -18.525 680.845 -18.195 ;
        RECT 679.155 -18.525 679.485 -18.195 ;
        RECT 677.795 -18.525 678.125 -18.195 ;
        RECT 675.075 -18.525 675.405 -18.195 ;
        RECT 673.715 -18.525 674.045 -18.195 ;
        RECT 672.355 -18.525 672.685 -18.195 ;
        RECT 670.995 -18.525 671.325 -18.195 ;
        RECT 669.635 -18.525 669.965 -18.195 ;
        RECT 668.275 -18.525 668.605 -18.195 ;
        RECT 666.915 -18.525 667.245 -18.195 ;
        RECT 665.555 -18.525 665.885 -18.195 ;
        RECT 664.195 -18.525 664.525 -18.195 ;
        RECT 662.835 -18.525 663.165 -18.195 ;
        RECT 660.115 -18.525 660.445 -18.195 ;
        RECT 658.755 -18.525 659.085 -18.195 ;
        RECT 657.395 -18.525 657.725 -18.195 ;
        RECT 656.035 -18.525 656.365 -18.195 ;
        RECT 654.675 -18.525 655.005 -18.195 ;
        RECT 653.315 -18.525 653.645 -18.195 ;
        RECT 815.155 -18.525 815.485 -18.195 ;
        RECT 813.795 -18.525 814.125 -18.195 ;
        RECT 812.435 -18.525 812.765 -18.195 ;
        RECT 808.355 -18.525 808.685 -18.195 ;
        RECT 806.995 -18.525 807.325 -18.195 ;
        RECT 805.635 -18.525 805.965 -18.195 ;
        RECT 804.275 -18.525 804.605 -18.195 ;
        RECT 802.915 -18.525 803.245 -18.195 ;
        RECT 801.555 -18.525 801.885 -18.195 ;
        RECT 800.195 -18.525 800.525 -18.195 ;
        RECT 798.835 -18.525 799.165 -18.195 ;
        RECT 797.475 -18.525 797.805 -18.195 ;
        RECT 793.395 -18.525 793.725 -18.195 ;
        RECT 792.035 -18.525 792.365 -18.195 ;
        RECT 790.675 -18.525 791.005 -18.195 ;
        RECT 789.315 -18.525 789.645 -18.195 ;
        RECT 787.955 -18.525 788.285 -18.195 ;
        RECT 786.595 -18.525 786.925 -18.195 ;
        RECT 785.235 -18.525 785.565 -18.195 ;
        RECT 783.875 -18.525 784.205 -18.195 ;
        RECT 782.515 -18.525 782.845 -18.195 ;
        RECT 778.435 -18.525 778.765 -18.195 ;
        RECT 777.405 -18.52 954.88 -18.2 ;
        RECT 953.875 -18.525 954.205 -18.195 ;
        RECT 952.515 -18.525 952.845 -18.195 ;
        RECT 951.155 -18.525 951.485 -18.195 ;
        RECT 949.795 -18.525 950.125 -18.195 ;
        RECT 948.435 -18.525 948.765 -18.195 ;
        RECT 947.075 -18.525 947.405 -18.195 ;
        RECT 945.715 -18.525 946.045 -18.195 ;
        RECT 944.355 -18.525 944.685 -18.195 ;
        RECT 942.995 -18.525 943.325 -18.195 ;
        RECT 941.635 -18.525 941.965 -18.195 ;
        RECT 940.275 -18.525 940.605 -18.195 ;
        RECT 938.915 -18.525 939.245 -18.195 ;
        RECT 937.555 -18.525 937.885 -18.195 ;
        RECT 936.195 -18.525 936.525 -18.195 ;
        RECT 934.835 -18.525 935.165 -18.195 ;
        RECT 933.475 -18.525 933.805 -18.195 ;
        RECT 932.115 -18.525 932.445 -18.195 ;
        RECT 930.755 -18.525 931.085 -18.195 ;
        RECT 928.035 -18.525 928.365 -18.195 ;
        RECT 926.675 -18.525 927.005 -18.195 ;
        RECT 925.315 -18.525 925.645 -18.195 ;
        RECT 923.955 -18.525 924.285 -18.195 ;
        RECT 922.595 -18.525 922.925 -18.195 ;
        RECT 921.235 -18.525 921.565 -18.195 ;
        RECT 919.875 -18.525 920.205 -18.195 ;
        RECT 918.515 -18.525 918.845 -18.195 ;
        RECT 917.155 -18.525 917.485 -18.195 ;
        RECT 913.075 -18.525 913.405 -18.195 ;
        RECT 911.715 -18.525 912.045 -18.195 ;
        RECT 910.355 -18.525 910.685 -18.195 ;
        RECT 908.995 -18.525 909.325 -18.195 ;
        RECT 907.635 -18.525 907.965 -18.195 ;
        RECT 906.275 -18.525 906.605 -18.195 ;
        RECT 904.915 -18.525 905.245 -18.195 ;
        RECT 903.555 -18.525 903.885 -18.195 ;
        RECT 902.195 -18.525 902.525 -18.195 ;
        RECT 898.115 -18.525 898.445 -18.195 ;
        RECT 896.755 -18.525 897.085 -18.195 ;
        RECT 895.395 -18.525 895.725 -18.195 ;
        RECT 894.035 -18.525 894.365 -18.195 ;
        RECT 892.675 -18.525 893.005 -18.195 ;
        RECT 891.315 -18.525 891.645 -18.195 ;
        RECT 889.955 -18.525 890.285 -18.195 ;
        RECT 888.595 -18.525 888.925 -18.195 ;
        RECT 887.235 -18.525 887.565 -18.195 ;
        RECT 883.155 -18.525 883.485 -18.195 ;
        RECT 881.795 -18.525 882.125 -18.195 ;
        RECT 880.435 -18.525 880.765 -18.195 ;
        RECT 879.075 -18.525 879.405 -18.195 ;
        RECT 877.715 -18.525 878.045 -18.195 ;
        RECT 876.355 -18.525 876.685 -18.195 ;
        RECT 874.995 -18.525 875.325 -18.195 ;
        RECT 873.635 -18.525 873.965 -18.195 ;
        RECT 872.275 -18.525 872.605 -18.195 ;
        RECT 868.195 -18.525 868.525 -18.195 ;
        RECT 866.835 -18.525 867.165 -18.195 ;
        RECT 865.475 -18.525 865.805 -18.195 ;
        RECT 864.115 -18.525 864.445 -18.195 ;
        RECT 862.755 -18.525 863.085 -18.195 ;
        RECT 861.395 -18.525 861.725 -18.195 ;
        RECT 860.035 -18.525 860.365 -18.195 ;
        RECT 858.675 -18.525 859.005 -18.195 ;
        RECT 857.315 -18.525 857.645 -18.195 ;
        RECT 853.235 -18.525 853.565 -18.195 ;
        RECT 851.875 -18.525 852.205 -18.195 ;
        RECT 850.515 -18.525 850.845 -18.195 ;
        RECT 849.155 -18.525 849.485 -18.195 ;
        RECT 847.795 -18.525 848.125 -18.195 ;
        RECT 846.435 -18.525 846.765 -18.195 ;
        RECT 845.075 -18.525 845.405 -18.195 ;
        RECT 843.715 -18.525 844.045 -18.195 ;
        RECT 842.355 -18.525 842.685 -18.195 ;
        RECT 838.275 -18.525 838.605 -18.195 ;
        RECT 836.915 -18.525 837.245 -18.195 ;
        RECT 835.555 -18.525 835.885 -18.195 ;
        RECT 834.195 -18.525 834.525 -18.195 ;
        RECT 832.835 -18.525 833.165 -18.195 ;
        RECT 831.475 -18.525 831.805 -18.195 ;
        RECT 830.115 -18.525 830.445 -18.195 ;
        RECT 828.755 -18.525 829.085 -18.195 ;
        RECT 827.395 -18.525 827.725 -18.195 ;
        RECT 823.315 -18.525 823.645 -18.195 ;
        RECT 821.955 -18.525 822.285 -18.195 ;
        RECT 820.595 -18.525 820.925 -18.195 ;
        RECT 819.235 -18.525 819.565 -18.195 ;
        RECT 817.875 -18.525 818.205 -18.195 ;
        RECT 816.515 -18.525 816.845 -18.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 -15.805 678.125 -15.475 ;
        RECT -1.52 -15.8 678.125 -15.48 ;
        RECT 676.435 -15.805 676.765 -15.475 ;
        RECT 675.075 -15.805 675.405 -15.475 ;
        RECT 673.715 -15.805 674.045 -15.475 ;
        RECT 672.355 -15.805 672.685 -15.475 ;
        RECT 670.995 -15.805 671.325 -15.475 ;
        RECT 669.635 -15.805 669.965 -15.475 ;
        RECT 668.275 -15.805 668.605 -15.475 ;
        RECT 666.915 -15.805 667.245 -15.475 ;
        RECT 665.555 -15.805 665.885 -15.475 ;
        RECT 664.195 -15.805 664.525 -15.475 ;
        RECT 662.835 -15.805 663.165 -15.475 ;
        RECT 661.475 -15.805 661.805 -15.475 ;
        RECT 660.115 -15.805 660.445 -15.475 ;
        RECT 658.755 -15.805 659.085 -15.475 ;
        RECT 657.395 -15.805 657.725 -15.475 ;
        RECT 656.035 -15.805 656.365 -15.475 ;
        RECT 654.675 -15.805 655.005 -15.475 ;
        RECT 653.315 -15.805 653.645 -15.475 ;
        RECT 651.955 -15.805 652.285 -15.475 ;
        RECT 650.595 -15.805 650.925 -15.475 ;
        RECT 649.235 -15.805 649.565 -15.475 ;
        RECT 647.875 -15.805 648.205 -15.475 ;
        RECT 646.515 -15.805 646.845 -15.475 ;
        RECT 645.155 -15.805 645.485 -15.475 ;
        RECT 643.795 -15.805 644.125 -15.475 ;
        RECT 642.435 -15.805 642.765 -15.475 ;
        RECT 641.075 -15.805 641.405 -15.475 ;
        RECT 639.715 -15.805 640.045 -15.475 ;
        RECT 638.355 -15.805 638.685 -15.475 ;
        RECT 636.995 -15.805 637.325 -15.475 ;
        RECT 635.635 -15.805 635.965 -15.475 ;
        RECT 634.275 -15.805 634.605 -15.475 ;
        RECT 632.915 -15.805 633.245 -15.475 ;
        RECT 631.555 -15.805 631.885 -15.475 ;
        RECT 630.195 -15.805 630.525 -15.475 ;
        RECT 628.835 -15.805 629.165 -15.475 ;
        RECT 627.475 -15.805 627.805 -15.475 ;
        RECT 626.115 -15.805 626.445 -15.475 ;
        RECT 624.755 -15.805 625.085 -15.475 ;
        RECT 623.395 -15.805 623.725 -15.475 ;
        RECT 622.035 -15.805 622.365 -15.475 ;
        RECT 620.675 -15.805 621.005 -15.475 ;
        RECT 619.315 -15.805 619.645 -15.475 ;
        RECT 617.955 -15.805 618.285 -15.475 ;
        RECT 616.595 -15.805 616.925 -15.475 ;
        RECT 615.235 -15.805 615.565 -15.475 ;
        RECT 613.875 -15.805 614.205 -15.475 ;
        RECT 612.515 -15.805 612.845 -15.475 ;
        RECT 611.155 -15.805 611.485 -15.475 ;
        RECT 609.795 -15.805 610.125 -15.475 ;
        RECT 608.435 -15.805 608.765 -15.475 ;
        RECT 607.075 -15.805 607.405 -15.475 ;
        RECT 605.715 -15.805 606.045 -15.475 ;
        RECT 604.355 -15.805 604.685 -15.475 ;
        RECT 602.995 -15.805 603.325 -15.475 ;
        RECT 601.635 -15.805 601.965 -15.475 ;
        RECT 600.275 -15.805 600.605 -15.475 ;
        RECT 598.915 -15.805 599.245 -15.475 ;
        RECT 597.555 -15.805 597.885 -15.475 ;
        RECT 596.195 -15.805 596.525 -15.475 ;
        RECT 594.835 -15.805 595.165 -15.475 ;
        RECT 593.475 -15.805 593.805 -15.475 ;
        RECT 592.115 -15.805 592.445 -15.475 ;
        RECT 590.755 -15.805 591.085 -15.475 ;
        RECT 589.395 -15.805 589.725 -15.475 ;
        RECT 588.035 -15.805 588.365 -15.475 ;
        RECT 586.675 -15.805 587.005 -15.475 ;
        RECT 585.315 -15.805 585.645 -15.475 ;
        RECT 583.955 -15.805 584.285 -15.475 ;
        RECT 582.595 -15.805 582.925 -15.475 ;
        RECT 581.235 -15.805 581.565 -15.475 ;
        RECT 579.875 -15.805 580.205 -15.475 ;
        RECT 578.515 -15.805 578.845 -15.475 ;
        RECT 577.155 -15.805 577.485 -15.475 ;
        RECT 575.795 -15.805 576.125 -15.475 ;
        RECT 574.435 -15.805 574.765 -15.475 ;
        RECT 573.075 -15.805 573.405 -15.475 ;
        RECT 571.715 -15.805 572.045 -15.475 ;
        RECT 570.355 -15.805 570.685 -15.475 ;
        RECT 568.995 -15.805 569.325 -15.475 ;
        RECT 567.635 -15.805 567.965 -15.475 ;
        RECT 566.275 -15.805 566.605 -15.475 ;
        RECT 564.915 -15.805 565.245 -15.475 ;
        RECT 563.555 -15.805 563.885 -15.475 ;
        RECT 562.195 -15.805 562.525 -15.475 ;
        RECT 560.835 -15.805 561.165 -15.475 ;
        RECT 559.475 -15.805 559.805 -15.475 ;
        RECT 558.115 -15.805 558.445 -15.475 ;
        RECT 556.755 -15.805 557.085 -15.475 ;
        RECT 555.395 -15.805 555.725 -15.475 ;
        RECT 554.035 -15.805 554.365 -15.475 ;
        RECT 552.675 -15.805 553.005 -15.475 ;
        RECT 551.315 -15.805 551.645 -15.475 ;
        RECT 549.955 -15.805 550.285 -15.475 ;
        RECT 548.595 -15.805 548.925 -15.475 ;
        RECT 547.235 -15.805 547.565 -15.475 ;
        RECT 545.875 -15.805 546.205 -15.475 ;
        RECT 544.515 -15.805 544.845 -15.475 ;
        RECT 543.155 -15.805 543.485 -15.475 ;
        RECT 541.795 -15.805 542.125 -15.475 ;
        RECT 540.435 -15.805 540.765 -15.475 ;
        RECT 539.075 -15.805 539.405 -15.475 ;
        RECT 537.715 -15.805 538.045 -15.475 ;
        RECT 536.355 -15.805 536.685 -15.475 ;
        RECT 534.995 -15.805 535.325 -15.475 ;
        RECT 533.635 -15.805 533.965 -15.475 ;
        RECT 532.275 -15.805 532.605 -15.475 ;
        RECT 530.915 -15.805 531.245 -15.475 ;
        RECT 529.555 -15.805 529.885 -15.475 ;
        RECT 528.195 -15.805 528.525 -15.475 ;
        RECT 526.835 -15.805 527.165 -15.475 ;
        RECT 525.475 -15.805 525.805 -15.475 ;
        RECT 524.115 -15.805 524.445 -15.475 ;
        RECT 522.755 -15.805 523.085 -15.475 ;
        RECT 521.395 -15.805 521.725 -15.475 ;
        RECT 520.035 -15.805 520.365 -15.475 ;
        RECT 518.675 -15.805 519.005 -15.475 ;
        RECT 517.315 -15.805 517.645 -15.475 ;
        RECT 515.955 -15.805 516.285 -15.475 ;
        RECT 514.595 -15.805 514.925 -15.475 ;
        RECT 513.235 -15.805 513.565 -15.475 ;
        RECT 511.875 -15.805 512.205 -15.475 ;
        RECT 510.515 -15.805 510.845 -15.475 ;
        RECT 509.155 -15.805 509.485 -15.475 ;
        RECT 507.795 -15.805 508.125 -15.475 ;
        RECT 506.435 -15.805 506.765 -15.475 ;
        RECT 505.075 -15.805 505.405 -15.475 ;
        RECT 503.715 -15.805 504.045 -15.475 ;
        RECT 502.355 -15.805 502.685 -15.475 ;
        RECT 500.995 -15.805 501.325 -15.475 ;
        RECT 499.635 -15.805 499.965 -15.475 ;
        RECT 498.275 -15.805 498.605 -15.475 ;
        RECT 496.915 -15.805 497.245 -15.475 ;
        RECT 495.555 -15.805 495.885 -15.475 ;
        RECT 494.195 -15.805 494.525 -15.475 ;
        RECT 492.835 -15.805 493.165 -15.475 ;
        RECT 491.475 -15.805 491.805 -15.475 ;
        RECT 490.115 -15.805 490.445 -15.475 ;
        RECT 488.755 -15.805 489.085 -15.475 ;
        RECT 487.395 -15.805 487.725 -15.475 ;
        RECT 486.035 -15.805 486.365 -15.475 ;
        RECT 484.675 -15.805 485.005 -15.475 ;
        RECT 483.315 -15.805 483.645 -15.475 ;
        RECT 481.955 -15.805 482.285 -15.475 ;
        RECT 480.595 -15.805 480.925 -15.475 ;
        RECT 479.235 -15.805 479.565 -15.475 ;
        RECT 477.875 -15.805 478.205 -15.475 ;
        RECT 476.515 -15.805 476.845 -15.475 ;
        RECT 475.155 -15.805 475.485 -15.475 ;
        RECT 473.795 -15.805 474.125 -15.475 ;
        RECT 472.435 -15.805 472.765 -15.475 ;
        RECT 471.075 -15.805 471.405 -15.475 ;
        RECT 469.715 -15.805 470.045 -15.475 ;
        RECT 468.355 -15.805 468.685 -15.475 ;
        RECT 466.995 -15.805 467.325 -15.475 ;
        RECT 465.635 -15.805 465.965 -15.475 ;
        RECT 464.275 -15.805 464.605 -15.475 ;
        RECT 462.915 -15.805 463.245 -15.475 ;
        RECT 461.555 -15.805 461.885 -15.475 ;
        RECT 460.195 -15.805 460.525 -15.475 ;
        RECT 458.835 -15.805 459.165 -15.475 ;
        RECT 457.475 -15.805 457.805 -15.475 ;
        RECT 456.115 -15.805 456.445 -15.475 ;
        RECT 454.755 -15.805 455.085 -15.475 ;
        RECT 453.395 -15.805 453.725 -15.475 ;
        RECT 452.035 -15.805 452.365 -15.475 ;
        RECT 450.675 -15.805 451.005 -15.475 ;
        RECT 449.315 -15.805 449.645 -15.475 ;
        RECT 447.955 -15.805 448.285 -15.475 ;
        RECT 446.595 -15.805 446.925 -15.475 ;
        RECT 445.235 -15.805 445.565 -15.475 ;
        RECT 443.875 -15.805 444.205 -15.475 ;
        RECT 442.515 -15.805 442.845 -15.475 ;
        RECT 441.155 -15.805 441.485 -15.475 ;
        RECT 439.795 -15.805 440.125 -15.475 ;
        RECT 438.435 -15.805 438.765 -15.475 ;
        RECT 437.075 -15.805 437.405 -15.475 ;
        RECT 435.715 -15.805 436.045 -15.475 ;
        RECT 434.355 -15.805 434.685 -15.475 ;
        RECT 432.995 -15.805 433.325 -15.475 ;
        RECT 431.635 -15.805 431.965 -15.475 ;
        RECT 430.275 -15.805 430.605 -15.475 ;
        RECT 428.915 -15.805 429.245 -15.475 ;
        RECT 427.555 -15.805 427.885 -15.475 ;
        RECT 426.195 -15.805 426.525 -15.475 ;
        RECT 424.835 -15.805 425.165 -15.475 ;
        RECT 423.475 -15.805 423.805 -15.475 ;
        RECT 422.115 -15.805 422.445 -15.475 ;
        RECT 420.755 -15.805 421.085 -15.475 ;
        RECT 419.395 -15.805 419.725 -15.475 ;
        RECT 418.035 -15.805 418.365 -15.475 ;
        RECT 416.675 -15.805 417.005 -15.475 ;
        RECT 415.315 -15.805 415.645 -15.475 ;
        RECT 413.955 -15.805 414.285 -15.475 ;
        RECT 412.595 -15.805 412.925 -15.475 ;
        RECT 411.235 -15.805 411.565 -15.475 ;
        RECT 409.875 -15.805 410.205 -15.475 ;
        RECT 408.515 -15.805 408.845 -15.475 ;
        RECT 407.155 -15.805 407.485 -15.475 ;
        RECT 405.795 -15.805 406.125 -15.475 ;
        RECT 404.435 -15.805 404.765 -15.475 ;
        RECT 403.075 -15.805 403.405 -15.475 ;
        RECT 401.715 -15.805 402.045 -15.475 ;
        RECT 400.355 -15.805 400.685 -15.475 ;
        RECT 398.995 -15.805 399.325 -15.475 ;
        RECT 397.635 -15.805 397.965 -15.475 ;
        RECT 396.275 -15.805 396.605 -15.475 ;
        RECT 394.915 -15.805 395.245 -15.475 ;
        RECT 393.555 -15.805 393.885 -15.475 ;
        RECT 392.195 -15.805 392.525 -15.475 ;
        RECT 390.835 -15.805 391.165 -15.475 ;
        RECT 389.475 -15.805 389.805 -15.475 ;
        RECT 388.115 -15.805 388.445 -15.475 ;
        RECT 386.755 -15.805 387.085 -15.475 ;
        RECT 385.395 -15.805 385.725 -15.475 ;
        RECT 384.035 -15.805 384.365 -15.475 ;
        RECT 382.675 -15.805 383.005 -15.475 ;
        RECT 381.315 -15.805 381.645 -15.475 ;
        RECT 379.955 -15.805 380.285 -15.475 ;
        RECT 378.595 -15.805 378.925 -15.475 ;
        RECT 377.235 -15.805 377.565 -15.475 ;
        RECT 375.875 -15.805 376.205 -15.475 ;
        RECT 374.515 -15.805 374.845 -15.475 ;
        RECT 373.155 -15.805 373.485 -15.475 ;
        RECT 371.795 -15.805 372.125 -15.475 ;
        RECT 370.435 -15.805 370.765 -15.475 ;
        RECT 369.075 -15.805 369.405 -15.475 ;
        RECT 367.715 -15.805 368.045 -15.475 ;
        RECT 366.355 -15.805 366.685 -15.475 ;
        RECT 364.995 -15.805 365.325 -15.475 ;
        RECT 363.635 -15.805 363.965 -15.475 ;
        RECT 362.275 -15.805 362.605 -15.475 ;
        RECT 360.915 -15.805 361.245 -15.475 ;
        RECT 359.555 -15.805 359.885 -15.475 ;
        RECT 358.195 -15.805 358.525 -15.475 ;
        RECT 356.835 -15.805 357.165 -15.475 ;
        RECT 355.475 -15.805 355.805 -15.475 ;
        RECT 354.115 -15.805 354.445 -15.475 ;
        RECT 352.755 -15.805 353.085 -15.475 ;
        RECT 351.395 -15.805 351.725 -15.475 ;
        RECT 350.035 -15.805 350.365 -15.475 ;
        RECT 348.675 -15.805 349.005 -15.475 ;
        RECT 347.315 -15.805 347.645 -15.475 ;
        RECT 345.955 -15.805 346.285 -15.475 ;
        RECT 344.595 -15.805 344.925 -15.475 ;
        RECT 343.235 -15.805 343.565 -15.475 ;
        RECT 341.875 -15.805 342.205 -15.475 ;
        RECT 340.515 -15.805 340.845 -15.475 ;
        RECT 339.155 -15.805 339.485 -15.475 ;
        RECT 337.795 -15.805 338.125 -15.475 ;
        RECT 336.435 -15.805 336.765 -15.475 ;
        RECT 335.075 -15.805 335.405 -15.475 ;
        RECT 333.715 -15.805 334.045 -15.475 ;
        RECT 332.355 -15.805 332.685 -15.475 ;
        RECT 330.995 -15.805 331.325 -15.475 ;
        RECT 329.635 -15.805 329.965 -15.475 ;
        RECT 328.275 -15.805 328.605 -15.475 ;
        RECT 326.915 -15.805 327.245 -15.475 ;
        RECT 325.555 -15.805 325.885 -15.475 ;
        RECT 324.195 -15.805 324.525 -15.475 ;
        RECT 322.835 -15.805 323.165 -15.475 ;
        RECT 321.475 -15.805 321.805 -15.475 ;
        RECT 320.115 -15.805 320.445 -15.475 ;
        RECT 318.755 -15.805 319.085 -15.475 ;
        RECT 317.395 -15.805 317.725 -15.475 ;
        RECT 316.035 -15.805 316.365 -15.475 ;
        RECT 314.675 -15.805 315.005 -15.475 ;
        RECT 313.315 -15.805 313.645 -15.475 ;
        RECT 311.955 -15.805 312.285 -15.475 ;
        RECT 310.595 -15.805 310.925 -15.475 ;
        RECT 309.235 -15.805 309.565 -15.475 ;
        RECT 307.875 -15.805 308.205 -15.475 ;
        RECT 306.515 -15.805 306.845 -15.475 ;
        RECT 305.155 -15.805 305.485 -15.475 ;
        RECT 303.795 -15.805 304.125 -15.475 ;
        RECT 302.435 -15.805 302.765 -15.475 ;
        RECT 301.075 -15.805 301.405 -15.475 ;
        RECT 299.715 -15.805 300.045 -15.475 ;
        RECT 298.355 -15.805 298.685 -15.475 ;
        RECT 296.995 -15.805 297.325 -15.475 ;
        RECT 295.635 -15.805 295.965 -15.475 ;
        RECT 294.275 -15.805 294.605 -15.475 ;
        RECT 292.915 -15.805 293.245 -15.475 ;
        RECT 291.555 -15.805 291.885 -15.475 ;
        RECT 290.195 -15.805 290.525 -15.475 ;
        RECT 288.835 -15.805 289.165 -15.475 ;
        RECT 287.475 -15.805 287.805 -15.475 ;
        RECT 286.115 -15.805 286.445 -15.475 ;
        RECT 284.755 -15.805 285.085 -15.475 ;
        RECT 283.395 -15.805 283.725 -15.475 ;
        RECT 282.035 -15.805 282.365 -15.475 ;
        RECT 280.675 -15.805 281.005 -15.475 ;
        RECT 279.315 -15.805 279.645 -15.475 ;
        RECT 277.955 -15.805 278.285 -15.475 ;
        RECT 276.595 -15.805 276.925 -15.475 ;
        RECT 275.235 -15.805 275.565 -15.475 ;
        RECT 273.875 -15.805 274.205 -15.475 ;
        RECT 272.515 -15.805 272.845 -15.475 ;
        RECT 271.155 -15.805 271.485 -15.475 ;
        RECT 269.795 -15.805 270.125 -15.475 ;
        RECT 268.435 -15.805 268.765 -15.475 ;
        RECT 267.075 -15.805 267.405 -15.475 ;
        RECT 265.715 -15.805 266.045 -15.475 ;
        RECT 264.355 -15.805 264.685 -15.475 ;
        RECT 262.995 -15.805 263.325 -15.475 ;
        RECT 261.635 -15.805 261.965 -15.475 ;
        RECT 260.275 -15.805 260.605 -15.475 ;
        RECT 258.915 -15.805 259.245 -15.475 ;
        RECT 257.555 -15.805 257.885 -15.475 ;
        RECT 256.195 -15.805 256.525 -15.475 ;
        RECT 254.835 -15.805 255.165 -15.475 ;
        RECT 253.475 -15.805 253.805 -15.475 ;
        RECT 252.115 -15.805 252.445 -15.475 ;
        RECT 250.755 -15.805 251.085 -15.475 ;
        RECT 249.395 -15.805 249.725 -15.475 ;
        RECT 248.035 -15.805 248.365 -15.475 ;
        RECT 246.675 -15.805 247.005 -15.475 ;
        RECT 245.315 -15.805 245.645 -15.475 ;
        RECT 243.955 -15.805 244.285 -15.475 ;
        RECT 242.595 -15.805 242.925 -15.475 ;
        RECT 241.235 -15.805 241.565 -15.475 ;
        RECT 239.875 -15.805 240.205 -15.475 ;
        RECT 238.515 -15.805 238.845 -15.475 ;
        RECT 237.155 -15.805 237.485 -15.475 ;
        RECT 235.795 -15.805 236.125 -15.475 ;
        RECT 234.435 -15.805 234.765 -15.475 ;
        RECT 233.075 -15.805 233.405 -15.475 ;
        RECT 231.715 -15.805 232.045 -15.475 ;
        RECT 230.355 -15.805 230.685 -15.475 ;
        RECT 228.995 -15.805 229.325 -15.475 ;
        RECT 227.635 -15.805 227.965 -15.475 ;
        RECT 226.275 -15.805 226.605 -15.475 ;
        RECT 224.915 -15.805 225.245 -15.475 ;
        RECT 223.555 -15.805 223.885 -15.475 ;
        RECT 222.195 -15.805 222.525 -15.475 ;
        RECT 220.835 -15.805 221.165 -15.475 ;
        RECT 219.475 -15.805 219.805 -15.475 ;
        RECT 218.115 -15.805 218.445 -15.475 ;
        RECT 216.755 -15.805 217.085 -15.475 ;
        RECT 215.395 -15.805 215.725 -15.475 ;
        RECT 214.035 -15.805 214.365 -15.475 ;
        RECT 212.675 -15.805 213.005 -15.475 ;
        RECT 211.315 -15.805 211.645 -15.475 ;
        RECT 209.955 -15.805 210.285 -15.475 ;
        RECT 208.595 -15.805 208.925 -15.475 ;
        RECT 207.235 -15.805 207.565 -15.475 ;
        RECT 205.875 -15.805 206.205 -15.475 ;
        RECT 204.515 -15.805 204.845 -15.475 ;
        RECT 203.155 -15.805 203.485 -15.475 ;
        RECT 201.795 -15.805 202.125 -15.475 ;
        RECT 200.435 -15.805 200.765 -15.475 ;
        RECT 199.075 -15.805 199.405 -15.475 ;
        RECT 197.715 -15.805 198.045 -15.475 ;
        RECT 196.355 -15.805 196.685 -15.475 ;
        RECT 194.995 -15.805 195.325 -15.475 ;
        RECT 193.635 -15.805 193.965 -15.475 ;
        RECT 192.275 -15.805 192.605 -15.475 ;
        RECT 190.915 -15.805 191.245 -15.475 ;
        RECT 189.555 -15.805 189.885 -15.475 ;
        RECT 188.195 -15.805 188.525 -15.475 ;
        RECT 186.835 -15.805 187.165 -15.475 ;
        RECT 185.475 -15.805 185.805 -15.475 ;
        RECT 184.115 -15.805 184.445 -15.475 ;
        RECT 182.755 -15.805 183.085 -15.475 ;
        RECT 181.395 -15.805 181.725 -15.475 ;
        RECT 180.035 -15.805 180.365 -15.475 ;
        RECT 178.675 -15.805 179.005 -15.475 ;
        RECT 177.315 -15.805 177.645 -15.475 ;
        RECT 175.955 -15.805 176.285 -15.475 ;
        RECT 174.595 -15.805 174.925 -15.475 ;
        RECT 173.235 -15.805 173.565 -15.475 ;
        RECT 171.875 -15.805 172.205 -15.475 ;
        RECT 170.515 -15.805 170.845 -15.475 ;
        RECT 169.155 -15.805 169.485 -15.475 ;
        RECT 167.795 -15.805 168.125 -15.475 ;
        RECT 166.435 -15.805 166.765 -15.475 ;
        RECT 165.075 -15.805 165.405 -15.475 ;
        RECT 163.715 -15.805 164.045 -15.475 ;
        RECT 162.355 -15.805 162.685 -15.475 ;
        RECT 160.995 -15.805 161.325 -15.475 ;
        RECT 159.635 -15.805 159.965 -15.475 ;
        RECT 158.275 -15.805 158.605 -15.475 ;
        RECT 156.915 -15.805 157.245 -15.475 ;
        RECT 155.555 -15.805 155.885 -15.475 ;
        RECT 154.195 -15.805 154.525 -15.475 ;
        RECT 152.835 -15.805 153.165 -15.475 ;
        RECT 151.475 -15.805 151.805 -15.475 ;
        RECT 150.115 -15.805 150.445 -15.475 ;
        RECT 148.755 -15.805 149.085 -15.475 ;
        RECT 147.395 -15.805 147.725 -15.475 ;
        RECT 146.035 -15.805 146.365 -15.475 ;
        RECT 144.675 -15.805 145.005 -15.475 ;
        RECT 143.315 -15.805 143.645 -15.475 ;
        RECT 141.955 -15.805 142.285 -15.475 ;
        RECT 140.595 -15.805 140.925 -15.475 ;
        RECT 139.235 -15.805 139.565 -15.475 ;
        RECT 137.875 -15.805 138.205 -15.475 ;
        RECT 136.515 -15.805 136.845 -15.475 ;
        RECT 135.155 -15.805 135.485 -15.475 ;
        RECT 133.795 -15.805 134.125 -15.475 ;
        RECT 132.435 -15.805 132.765 -15.475 ;
        RECT 131.075 -15.805 131.405 -15.475 ;
        RECT 129.715 -15.805 130.045 -15.475 ;
        RECT 128.355 -15.805 128.685 -15.475 ;
        RECT 126.995 -15.805 127.325 -15.475 ;
        RECT 125.635 -15.805 125.965 -15.475 ;
        RECT 124.275 -15.805 124.605 -15.475 ;
        RECT 122.915 -15.805 123.245 -15.475 ;
        RECT 121.555 -15.805 121.885 -15.475 ;
        RECT 120.195 -15.805 120.525 -15.475 ;
        RECT 118.835 -15.805 119.165 -15.475 ;
        RECT 117.475 -15.805 117.805 -15.475 ;
        RECT 116.115 -15.805 116.445 -15.475 ;
        RECT 114.755 -15.805 115.085 -15.475 ;
        RECT 113.395 -15.805 113.725 -15.475 ;
        RECT 112.035 -15.805 112.365 -15.475 ;
        RECT 110.675 -15.805 111.005 -15.475 ;
        RECT 109.315 -15.805 109.645 -15.475 ;
        RECT 107.955 -15.805 108.285 -15.475 ;
        RECT 106.595 -15.805 106.925 -15.475 ;
        RECT 105.235 -15.805 105.565 -15.475 ;
        RECT 103.875 -15.805 104.205 -15.475 ;
        RECT 102.515 -15.805 102.845 -15.475 ;
        RECT 101.155 -15.805 101.485 -15.475 ;
        RECT 99.795 -15.805 100.125 -15.475 ;
        RECT 98.435 -15.805 98.765 -15.475 ;
        RECT 97.075 -15.805 97.405 -15.475 ;
        RECT 95.715 -15.805 96.045 -15.475 ;
        RECT 94.355 -15.805 94.685 -15.475 ;
        RECT 92.995 -15.805 93.325 -15.475 ;
        RECT 91.635 -15.805 91.965 -15.475 ;
        RECT 90.275 -15.805 90.605 -15.475 ;
        RECT 88.915 -15.805 89.245 -15.475 ;
        RECT 87.555 -15.805 87.885 -15.475 ;
        RECT 86.195 -15.805 86.525 -15.475 ;
        RECT 84.835 -15.805 85.165 -15.475 ;
        RECT 83.475 -15.805 83.805 -15.475 ;
        RECT 82.115 -15.805 82.445 -15.475 ;
        RECT 80.755 -15.805 81.085 -15.475 ;
        RECT 79.395 -15.805 79.725 -15.475 ;
        RECT 78.035 -15.805 78.365 -15.475 ;
        RECT 76.675 -15.805 77.005 -15.475 ;
        RECT 75.315 -15.805 75.645 -15.475 ;
        RECT 73.955 -15.805 74.285 -15.475 ;
        RECT 72.595 -15.805 72.925 -15.475 ;
        RECT 71.235 -15.805 71.565 -15.475 ;
        RECT 69.875 -15.805 70.205 -15.475 ;
        RECT 68.515 -15.805 68.845 -15.475 ;
        RECT 67.155 -15.805 67.485 -15.475 ;
        RECT 65.795 -15.805 66.125 -15.475 ;
        RECT 64.435 -15.805 64.765 -15.475 ;
        RECT 63.075 -15.805 63.405 -15.475 ;
        RECT 61.715 -15.805 62.045 -15.475 ;
        RECT 60.355 -15.805 60.685 -15.475 ;
        RECT 58.995 -15.805 59.325 -15.475 ;
        RECT 57.635 -15.805 57.965 -15.475 ;
        RECT 56.275 -15.805 56.605 -15.475 ;
        RECT 54.915 -15.805 55.245 -15.475 ;
        RECT 53.555 -15.805 53.885 -15.475 ;
        RECT 52.195 -15.805 52.525 -15.475 ;
        RECT 50.835 -15.805 51.165 -15.475 ;
        RECT 49.475 -15.805 49.805 -15.475 ;
        RECT 48.115 -15.805 48.445 -15.475 ;
        RECT 46.755 -15.805 47.085 -15.475 ;
        RECT 45.395 -15.805 45.725 -15.475 ;
        RECT 44.035 -15.805 44.365 -15.475 ;
        RECT 42.675 -15.805 43.005 -15.475 ;
        RECT 41.315 -15.805 41.645 -15.475 ;
        RECT 39.955 -15.805 40.285 -15.475 ;
        RECT 38.595 -15.805 38.925 -15.475 ;
        RECT 37.235 -15.805 37.565 -15.475 ;
        RECT 35.875 -15.805 36.205 -15.475 ;
        RECT 34.515 -15.805 34.845 -15.475 ;
        RECT 33.155 -15.805 33.485 -15.475 ;
        RECT 31.795 -15.805 32.125 -15.475 ;
        RECT 30.435 -15.805 30.765 -15.475 ;
        RECT 29.075 -15.805 29.405 -15.475 ;
        RECT 27.715 -15.805 28.045 -15.475 ;
        RECT 26.355 -15.805 26.685 -15.475 ;
        RECT 24.995 -15.805 25.325 -15.475 ;
        RECT 23.635 -15.805 23.965 -15.475 ;
        RECT 22.275 -15.805 22.605 -15.475 ;
        RECT 20.915 -15.805 21.245 -15.475 ;
        RECT 19.555 -15.805 19.885 -15.475 ;
        RECT 18.195 -15.805 18.525 -15.475 ;
        RECT 16.835 -15.805 17.165 -15.475 ;
        RECT 15.475 -15.805 15.805 -15.475 ;
        RECT 14.115 -15.805 14.445 -15.475 ;
        RECT 12.755 -15.805 13.085 -15.475 ;
        RECT 11.395 -15.805 11.725 -15.475 ;
        RECT 10.035 -15.805 10.365 -15.475 ;
        RECT 8.675 -15.805 9.005 -15.475 ;
        RECT 7.315 -15.805 7.645 -15.475 ;
        RECT 5.955 -15.805 6.285 -15.475 ;
        RECT 4.595 -15.805 4.925 -15.475 ;
        RECT 3.235 -15.805 3.565 -15.475 ;
        RECT 1.875 -15.805 2.205 -15.475 ;
        RECT 0.515 -15.805 0.845 -15.475 ;
        RECT -0.845 -15.805 -0.515 -15.475 ;
        RECT 678.125 -15.8 954.88 -15.48 ;
        RECT 953.875 -15.805 954.205 -15.475 ;
        RECT 952.515 -15.805 952.845 -15.475 ;
        RECT 951.155 -15.805 951.485 -15.475 ;
        RECT 949.795 -15.805 950.125 -15.475 ;
        RECT 948.435 -15.805 948.765 -15.475 ;
        RECT 947.075 -15.805 947.405 -15.475 ;
        RECT 945.715 -15.805 946.045 -15.475 ;
        RECT 944.355 -15.805 944.685 -15.475 ;
        RECT 942.995 -15.805 943.325 -15.475 ;
        RECT 941.635 -15.805 941.965 -15.475 ;
        RECT 940.275 -15.805 940.605 -15.475 ;
        RECT 938.915 -15.805 939.245 -15.475 ;
        RECT 937.555 -15.805 937.885 -15.475 ;
        RECT 936.195 -15.805 936.525 -15.475 ;
        RECT 934.835 -15.805 935.165 -15.475 ;
        RECT 933.475 -15.805 933.805 -15.475 ;
        RECT 932.115 -15.805 932.445 -15.475 ;
        RECT 930.755 -15.805 931.085 -15.475 ;
        RECT 929.395 -15.805 929.725 -15.475 ;
        RECT 928.035 -15.805 928.365 -15.475 ;
        RECT 926.675 -15.805 927.005 -15.475 ;
        RECT 925.315 -15.805 925.645 -15.475 ;
        RECT 923.955 -15.805 924.285 -15.475 ;
        RECT 922.595 -15.805 922.925 -15.475 ;
        RECT 921.235 -15.805 921.565 -15.475 ;
        RECT 919.875 -15.805 920.205 -15.475 ;
        RECT 918.515 -15.805 918.845 -15.475 ;
        RECT 917.155 -15.805 917.485 -15.475 ;
        RECT 915.795 -15.805 916.125 -15.475 ;
        RECT 914.435 -15.805 914.765 -15.475 ;
        RECT 913.075 -15.805 913.405 -15.475 ;
        RECT 911.715 -15.805 912.045 -15.475 ;
        RECT 910.355 -15.805 910.685 -15.475 ;
        RECT 908.995 -15.805 909.325 -15.475 ;
        RECT 907.635 -15.805 907.965 -15.475 ;
        RECT 906.275 -15.805 906.605 -15.475 ;
        RECT 904.915 -15.805 905.245 -15.475 ;
        RECT 903.555 -15.805 903.885 -15.475 ;
        RECT 902.195 -15.805 902.525 -15.475 ;
        RECT 900.835 -15.805 901.165 -15.475 ;
        RECT 899.475 -15.805 899.805 -15.475 ;
        RECT 898.115 -15.805 898.445 -15.475 ;
        RECT 896.755 -15.805 897.085 -15.475 ;
        RECT 895.395 -15.805 895.725 -15.475 ;
        RECT 894.035 -15.805 894.365 -15.475 ;
        RECT 892.675 -15.805 893.005 -15.475 ;
        RECT 891.315 -15.805 891.645 -15.475 ;
        RECT 889.955 -15.805 890.285 -15.475 ;
        RECT 888.595 -15.805 888.925 -15.475 ;
        RECT 887.235 -15.805 887.565 -15.475 ;
        RECT 885.875 -15.805 886.205 -15.475 ;
        RECT 884.515 -15.805 884.845 -15.475 ;
        RECT 883.155 -15.805 883.485 -15.475 ;
        RECT 881.795 -15.805 882.125 -15.475 ;
        RECT 880.435 -15.805 880.765 -15.475 ;
        RECT 879.075 -15.805 879.405 -15.475 ;
        RECT 877.715 -15.805 878.045 -15.475 ;
        RECT 876.355 -15.805 876.685 -15.475 ;
        RECT 874.995 -15.805 875.325 -15.475 ;
        RECT 873.635 -15.805 873.965 -15.475 ;
        RECT 872.275 -15.805 872.605 -15.475 ;
        RECT 870.915 -15.805 871.245 -15.475 ;
        RECT 869.555 -15.805 869.885 -15.475 ;
        RECT 868.195 -15.805 868.525 -15.475 ;
        RECT 866.835 -15.805 867.165 -15.475 ;
        RECT 865.475 -15.805 865.805 -15.475 ;
        RECT 864.115 -15.805 864.445 -15.475 ;
        RECT 862.755 -15.805 863.085 -15.475 ;
        RECT 861.395 -15.805 861.725 -15.475 ;
        RECT 860.035 -15.805 860.365 -15.475 ;
        RECT 858.675 -15.805 859.005 -15.475 ;
        RECT 857.315 -15.805 857.645 -15.475 ;
        RECT 855.955 -15.805 856.285 -15.475 ;
        RECT 854.595 -15.805 854.925 -15.475 ;
        RECT 853.235 -15.805 853.565 -15.475 ;
        RECT 851.875 -15.805 852.205 -15.475 ;
        RECT 850.515 -15.805 850.845 -15.475 ;
        RECT 849.155 -15.805 849.485 -15.475 ;
        RECT 847.795 -15.805 848.125 -15.475 ;
        RECT 846.435 -15.805 846.765 -15.475 ;
        RECT 845.075 -15.805 845.405 -15.475 ;
        RECT 843.715 -15.805 844.045 -15.475 ;
        RECT 842.355 -15.805 842.685 -15.475 ;
        RECT 840.995 -15.805 841.325 -15.475 ;
        RECT 839.635 -15.805 839.965 -15.475 ;
        RECT 838.275 -15.805 838.605 -15.475 ;
        RECT 836.915 -15.805 837.245 -15.475 ;
        RECT 835.555 -15.805 835.885 -15.475 ;
        RECT 834.195 -15.805 834.525 -15.475 ;
        RECT 832.835 -15.805 833.165 -15.475 ;
        RECT 831.475 -15.805 831.805 -15.475 ;
        RECT 830.115 -15.805 830.445 -15.475 ;
        RECT 828.755 -15.805 829.085 -15.475 ;
        RECT 827.395 -15.805 827.725 -15.475 ;
        RECT 826.035 -15.805 826.365 -15.475 ;
        RECT 824.675 -15.805 825.005 -15.475 ;
        RECT 823.315 -15.805 823.645 -15.475 ;
        RECT 821.955 -15.805 822.285 -15.475 ;
        RECT 820.595 -15.805 820.925 -15.475 ;
        RECT 819.235 -15.805 819.565 -15.475 ;
        RECT 817.875 -15.805 818.205 -15.475 ;
        RECT 816.515 -15.805 816.845 -15.475 ;
        RECT 815.155 -15.805 815.485 -15.475 ;
        RECT 813.795 -15.805 814.125 -15.475 ;
        RECT 812.435 -15.805 812.765 -15.475 ;
        RECT 811.075 -15.805 811.405 -15.475 ;
        RECT 809.715 -15.805 810.045 -15.475 ;
        RECT 808.355 -15.805 808.685 -15.475 ;
        RECT 806.995 -15.805 807.325 -15.475 ;
        RECT 805.635 -15.805 805.965 -15.475 ;
        RECT 804.275 -15.805 804.605 -15.475 ;
        RECT 802.915 -15.805 803.245 -15.475 ;
        RECT 801.555 -15.805 801.885 -15.475 ;
        RECT 800.195 -15.805 800.525 -15.475 ;
        RECT 798.835 -15.805 799.165 -15.475 ;
        RECT 797.475 -15.805 797.805 -15.475 ;
        RECT 796.115 -15.805 796.445 -15.475 ;
        RECT 794.755 -15.805 795.085 -15.475 ;
        RECT 793.395 -15.805 793.725 -15.475 ;
        RECT 792.035 -15.805 792.365 -15.475 ;
        RECT 790.675 -15.805 791.005 -15.475 ;
        RECT 789.315 -15.805 789.645 -15.475 ;
        RECT 787.955 -15.805 788.285 -15.475 ;
        RECT 786.595 -15.805 786.925 -15.475 ;
        RECT 785.235 -15.805 785.565 -15.475 ;
        RECT 783.875 -15.805 784.205 -15.475 ;
        RECT 782.515 -15.805 782.845 -15.475 ;
        RECT 781.155 -15.805 781.485 -15.475 ;
        RECT 779.795 -15.805 780.125 -15.475 ;
        RECT 778.435 -15.805 778.765 -15.475 ;
        RECT 777.075 -15.805 777.405 -15.475 ;
        RECT 775.715 -15.805 776.045 -15.475 ;
        RECT 774.355 -15.805 774.685 -15.475 ;
        RECT 772.995 -15.805 773.325 -15.475 ;
        RECT 771.635 -15.805 771.965 -15.475 ;
        RECT 770.275 -15.805 770.605 -15.475 ;
        RECT 768.915 -15.805 769.245 -15.475 ;
        RECT 767.555 -15.805 767.885 -15.475 ;
        RECT 766.195 -15.805 766.525 -15.475 ;
        RECT 764.835 -15.805 765.165 -15.475 ;
        RECT 763.475 -15.805 763.805 -15.475 ;
        RECT 762.115 -15.805 762.445 -15.475 ;
        RECT 760.755 -15.805 761.085 -15.475 ;
        RECT 759.395 -15.805 759.725 -15.475 ;
        RECT 758.035 -15.805 758.365 -15.475 ;
        RECT 756.675 -15.805 757.005 -15.475 ;
        RECT 755.315 -15.805 755.645 -15.475 ;
        RECT 753.955 -15.805 754.285 -15.475 ;
        RECT 752.595 -15.805 752.925 -15.475 ;
        RECT 751.235 -15.805 751.565 -15.475 ;
        RECT 749.875 -15.805 750.205 -15.475 ;
        RECT 748.515 -15.805 748.845 -15.475 ;
        RECT 747.155 -15.805 747.485 -15.475 ;
        RECT 745.795 -15.805 746.125 -15.475 ;
        RECT 744.435 -15.805 744.765 -15.475 ;
        RECT 743.075 -15.805 743.405 -15.475 ;
        RECT 741.715 -15.805 742.045 -15.475 ;
        RECT 740.355 -15.805 740.685 -15.475 ;
        RECT 738.995 -15.805 739.325 -15.475 ;
        RECT 737.635 -15.805 737.965 -15.475 ;
        RECT 736.275 -15.805 736.605 -15.475 ;
        RECT 734.915 -15.805 735.245 -15.475 ;
        RECT 733.555 -15.805 733.885 -15.475 ;
        RECT 732.195 -15.805 732.525 -15.475 ;
        RECT 730.835 -15.805 731.165 -15.475 ;
        RECT 729.475 -15.805 729.805 -15.475 ;
        RECT 728.115 -15.805 728.445 -15.475 ;
        RECT 726.755 -15.805 727.085 -15.475 ;
        RECT 725.395 -15.805 725.725 -15.475 ;
        RECT 724.035 -15.805 724.365 -15.475 ;
        RECT 722.675 -15.805 723.005 -15.475 ;
        RECT 721.315 -15.805 721.645 -15.475 ;
        RECT 719.955 -15.805 720.285 -15.475 ;
        RECT 718.595 -15.805 718.925 -15.475 ;
        RECT 717.235 -15.805 717.565 -15.475 ;
        RECT 715.875 -15.805 716.205 -15.475 ;
        RECT 714.515 -15.805 714.845 -15.475 ;
        RECT 713.155 -15.805 713.485 -15.475 ;
        RECT 711.795 -15.805 712.125 -15.475 ;
        RECT 710.435 -15.805 710.765 -15.475 ;
        RECT 709.075 -15.805 709.405 -15.475 ;
        RECT 707.715 -15.805 708.045 -15.475 ;
        RECT 706.355 -15.805 706.685 -15.475 ;
        RECT 704.995 -15.805 705.325 -15.475 ;
        RECT 703.635 -15.805 703.965 -15.475 ;
        RECT 702.275 -15.805 702.605 -15.475 ;
        RECT 700.915 -15.805 701.245 -15.475 ;
        RECT 699.555 -15.805 699.885 -15.475 ;
        RECT 698.195 -15.805 698.525 -15.475 ;
        RECT 696.835 -15.805 697.165 -15.475 ;
        RECT 695.475 -15.805 695.805 -15.475 ;
        RECT 694.115 -15.805 694.445 -15.475 ;
        RECT 692.755 -15.805 693.085 -15.475 ;
        RECT 691.395 -15.805 691.725 -15.475 ;
        RECT 690.035 -15.805 690.365 -15.475 ;
        RECT 688.675 -15.805 689.005 -15.475 ;
        RECT 687.315 -15.805 687.645 -15.475 ;
        RECT 685.955 -15.805 686.285 -15.475 ;
        RECT 684.595 -15.805 684.925 -15.475 ;
        RECT 683.235 -15.805 683.565 -15.475 ;
        RECT 681.875 -15.805 682.205 -15.475 ;
        RECT 680.515 -15.805 680.845 -15.475 ;
        RECT 679.155 -15.805 679.485 -15.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -17.165 123.245 -16.835 ;
        RECT 121.555 -17.165 121.885 -16.835 ;
        RECT 120.195 -17.165 120.525 -16.835 ;
        RECT 118.835 -17.165 119.165 -16.835 ;
        RECT 117.475 -17.165 117.805 -16.835 ;
        RECT 116.115 -17.165 116.445 -16.835 ;
        RECT 114.755 -17.165 115.085 -16.835 ;
        RECT 113.395 -17.165 113.725 -16.835 ;
        RECT 112.035 -17.165 112.365 -16.835 ;
        RECT 110.675 -17.165 111.005 -16.835 ;
        RECT 109.315 -17.165 109.645 -16.835 ;
        RECT 107.955 -17.165 108.285 -16.835 ;
        RECT 106.595 -17.165 106.925 -16.835 ;
        RECT 105.235 -17.165 105.565 -16.835 ;
        RECT 103.875 -17.165 104.205 -16.835 ;
        RECT 102.515 -17.165 102.845 -16.835 ;
        RECT 101.155 -17.165 101.485 -16.835 ;
        RECT 99.795 -17.165 100.125 -16.835 ;
        RECT 98.435 -17.165 98.765 -16.835 ;
        RECT 97.075 -17.165 97.405 -16.835 ;
        RECT 95.715 -17.165 96.045 -16.835 ;
        RECT 94.355 -17.165 94.685 -16.835 ;
        RECT 92.995 -17.165 93.325 -16.835 ;
        RECT 91.635 -17.165 91.965 -16.835 ;
        RECT 90.275 -17.165 90.605 -16.835 ;
        RECT 88.915 -17.165 89.245 -16.835 ;
        RECT 87.555 -17.165 87.885 -16.835 ;
        RECT 86.195 -17.165 86.525 -16.835 ;
        RECT 84.835 -17.165 85.165 -16.835 ;
        RECT 83.475 -17.165 83.805 -16.835 ;
        RECT 82.115 -17.165 82.445 -16.835 ;
        RECT 80.755 -17.165 81.085 -16.835 ;
        RECT 79.395 -17.165 79.725 -16.835 ;
        RECT 78.035 -17.165 78.365 -16.835 ;
        RECT 76.675 -17.165 77.005 -16.835 ;
        RECT 75.315 -17.165 75.645 -16.835 ;
        RECT 73.955 -17.165 74.285 -16.835 ;
        RECT 72.595 -17.165 72.925 -16.835 ;
        RECT 71.235 -17.165 71.565 -16.835 ;
        RECT 69.875 -17.165 70.205 -16.835 ;
        RECT 68.515 -17.165 68.845 -16.835 ;
        RECT 67.155 -17.165 67.485 -16.835 ;
        RECT 65.795 -17.165 66.125 -16.835 ;
        RECT 64.435 -17.165 64.765 -16.835 ;
        RECT 63.075 -17.165 63.405 -16.835 ;
        RECT 61.715 -17.165 62.045 -16.835 ;
        RECT 60.355 -17.165 60.685 -16.835 ;
        RECT 58.995 -17.165 59.325 -16.835 ;
        RECT 57.635 -17.165 57.965 -16.835 ;
        RECT 56.275 -17.165 56.605 -16.835 ;
        RECT 54.915 -17.165 55.245 -16.835 ;
        RECT 53.555 -17.165 53.885 -16.835 ;
        RECT 52.195 -17.165 52.525 -16.835 ;
        RECT 50.835 -17.165 51.165 -16.835 ;
        RECT 49.475 -17.165 49.805 -16.835 ;
        RECT 48.115 -17.165 48.445 -16.835 ;
        RECT 46.755 -17.165 47.085 -16.835 ;
        RECT 45.395 -17.165 45.725 -16.835 ;
        RECT 44.035 -17.165 44.365 -16.835 ;
        RECT 42.675 -17.165 43.005 -16.835 ;
        RECT 41.315 -17.165 41.645 -16.835 ;
        RECT 39.955 -17.165 40.285 -16.835 ;
        RECT 38.595 -17.165 38.925 -16.835 ;
        RECT 37.235 -17.165 37.565 -16.835 ;
        RECT 35.875 -17.165 36.205 -16.835 ;
        RECT 34.515 -17.165 34.845 -16.835 ;
        RECT 33.155 -17.165 33.485 -16.835 ;
        RECT 31.795 -17.165 32.125 -16.835 ;
        RECT 30.435 -17.165 30.765 -16.835 ;
        RECT 29.075 -17.165 29.405 -16.835 ;
        RECT 27.715 -17.165 28.045 -16.835 ;
        RECT 26.355 -17.165 26.685 -16.835 ;
        RECT 24.995 -17.165 25.325 -16.835 ;
        RECT 23.635 -17.165 23.965 -16.835 ;
        RECT 22.275 -17.165 22.605 -16.835 ;
        RECT 20.915 -17.165 21.245 -16.835 ;
        RECT 19.555 -17.165 19.885 -16.835 ;
        RECT 18.195 -17.165 18.525 -16.835 ;
        RECT 16.835 -17.165 17.165 -16.835 ;
        RECT 15.475 -17.165 15.805 -16.835 ;
        RECT 14.115 -17.165 14.445 -16.835 ;
        RECT 12.755 -17.165 13.085 -16.835 ;
        RECT 11.395 -17.165 11.725 -16.835 ;
        RECT 10.035 -17.165 10.365 -16.835 ;
        RECT 8.675 -17.165 9.005 -16.835 ;
        RECT 7.315 -17.165 7.645 -16.835 ;
        RECT 5.955 -17.165 6.285 -16.835 ;
        RECT 4.595 -17.165 4.925 -16.835 ;
        RECT 3.235 -17.165 3.565 -16.835 ;
        RECT 1.875 -17.165 2.205 -16.835 ;
        RECT 0.515 -17.165 0.845 -16.835 ;
        RECT -0.845 -17.165 -0.515 -16.835 ;
        RECT 677.795 -17.165 678.125 -16.835 ;
        RECT -1.52 -17.16 678.125 -16.84 ;
        RECT 676.435 -17.165 676.765 -16.835 ;
        RECT 675.075 -17.165 675.405 -16.835 ;
        RECT 673.715 -17.165 674.045 -16.835 ;
        RECT 672.355 -17.165 672.685 -16.835 ;
        RECT 670.995 -17.165 671.325 -16.835 ;
        RECT 669.635 -17.165 669.965 -16.835 ;
        RECT 668.275 -17.165 668.605 -16.835 ;
        RECT 666.915 -17.165 667.245 -16.835 ;
        RECT 665.555 -17.165 665.885 -16.835 ;
        RECT 664.195 -17.165 664.525 -16.835 ;
        RECT 662.835 -17.165 663.165 -16.835 ;
        RECT 661.475 -17.165 661.805 -16.835 ;
        RECT 660.115 -17.165 660.445 -16.835 ;
        RECT 658.755 -17.165 659.085 -16.835 ;
        RECT 657.395 -17.165 657.725 -16.835 ;
        RECT 656.035 -17.165 656.365 -16.835 ;
        RECT 654.675 -17.165 655.005 -16.835 ;
        RECT 653.315 -17.165 653.645 -16.835 ;
        RECT 651.955 -17.165 652.285 -16.835 ;
        RECT 650.595 -17.165 650.925 -16.835 ;
        RECT 649.235 -17.165 649.565 -16.835 ;
        RECT 647.875 -17.165 648.205 -16.835 ;
        RECT 646.515 -17.165 646.845 -16.835 ;
        RECT 645.155 -17.165 645.485 -16.835 ;
        RECT 643.795 -17.165 644.125 -16.835 ;
        RECT 642.435 -17.165 642.765 -16.835 ;
        RECT 641.075 -17.165 641.405 -16.835 ;
        RECT 639.715 -17.165 640.045 -16.835 ;
        RECT 638.355 -17.165 638.685 -16.835 ;
        RECT 636.995 -17.165 637.325 -16.835 ;
        RECT 635.635 -17.165 635.965 -16.835 ;
        RECT 634.275 -17.165 634.605 -16.835 ;
        RECT 632.915 -17.165 633.245 -16.835 ;
        RECT 631.555 -17.165 631.885 -16.835 ;
        RECT 630.195 -17.165 630.525 -16.835 ;
        RECT 628.835 -17.165 629.165 -16.835 ;
        RECT 627.475 -17.165 627.805 -16.835 ;
        RECT 626.115 -17.165 626.445 -16.835 ;
        RECT 624.755 -17.165 625.085 -16.835 ;
        RECT 623.395 -17.165 623.725 -16.835 ;
        RECT 622.035 -17.165 622.365 -16.835 ;
        RECT 620.675 -17.165 621.005 -16.835 ;
        RECT 619.315 -17.165 619.645 -16.835 ;
        RECT 617.955 -17.165 618.285 -16.835 ;
        RECT 616.595 -17.165 616.925 -16.835 ;
        RECT 615.235 -17.165 615.565 -16.835 ;
        RECT 613.875 -17.165 614.205 -16.835 ;
        RECT 612.515 -17.165 612.845 -16.835 ;
        RECT 611.155 -17.165 611.485 -16.835 ;
        RECT 609.795 -17.165 610.125 -16.835 ;
        RECT 608.435 -17.165 608.765 -16.835 ;
        RECT 607.075 -17.165 607.405 -16.835 ;
        RECT 605.715 -17.165 606.045 -16.835 ;
        RECT 604.355 -17.165 604.685 -16.835 ;
        RECT 602.995 -17.165 603.325 -16.835 ;
        RECT 601.635 -17.165 601.965 -16.835 ;
        RECT 600.275 -17.165 600.605 -16.835 ;
        RECT 598.915 -17.165 599.245 -16.835 ;
        RECT 597.555 -17.165 597.885 -16.835 ;
        RECT 596.195 -17.165 596.525 -16.835 ;
        RECT 594.835 -17.165 595.165 -16.835 ;
        RECT 593.475 -17.165 593.805 -16.835 ;
        RECT 592.115 -17.165 592.445 -16.835 ;
        RECT 590.755 -17.165 591.085 -16.835 ;
        RECT 589.395 -17.165 589.725 -16.835 ;
        RECT 588.035 -17.165 588.365 -16.835 ;
        RECT 586.675 -17.165 587.005 -16.835 ;
        RECT 585.315 -17.165 585.645 -16.835 ;
        RECT 583.955 -17.165 584.285 -16.835 ;
        RECT 582.595 -17.165 582.925 -16.835 ;
        RECT 581.235 -17.165 581.565 -16.835 ;
        RECT 579.875 -17.165 580.205 -16.835 ;
        RECT 578.515 -17.165 578.845 -16.835 ;
        RECT 577.155 -17.165 577.485 -16.835 ;
        RECT 575.795 -17.165 576.125 -16.835 ;
        RECT 574.435 -17.165 574.765 -16.835 ;
        RECT 573.075 -17.165 573.405 -16.835 ;
        RECT 571.715 -17.165 572.045 -16.835 ;
        RECT 570.355 -17.165 570.685 -16.835 ;
        RECT 568.995 -17.165 569.325 -16.835 ;
        RECT 567.635 -17.165 567.965 -16.835 ;
        RECT 566.275 -17.165 566.605 -16.835 ;
        RECT 564.915 -17.165 565.245 -16.835 ;
        RECT 563.555 -17.165 563.885 -16.835 ;
        RECT 562.195 -17.165 562.525 -16.835 ;
        RECT 560.835 -17.165 561.165 -16.835 ;
        RECT 559.475 -17.165 559.805 -16.835 ;
        RECT 558.115 -17.165 558.445 -16.835 ;
        RECT 556.755 -17.165 557.085 -16.835 ;
        RECT 555.395 -17.165 555.725 -16.835 ;
        RECT 554.035 -17.165 554.365 -16.835 ;
        RECT 552.675 -17.165 553.005 -16.835 ;
        RECT 551.315 -17.165 551.645 -16.835 ;
        RECT 549.955 -17.165 550.285 -16.835 ;
        RECT 548.595 -17.165 548.925 -16.835 ;
        RECT 547.235 -17.165 547.565 -16.835 ;
        RECT 545.875 -17.165 546.205 -16.835 ;
        RECT 544.515 -17.165 544.845 -16.835 ;
        RECT 543.155 -17.165 543.485 -16.835 ;
        RECT 541.795 -17.165 542.125 -16.835 ;
        RECT 540.435 -17.165 540.765 -16.835 ;
        RECT 539.075 -17.165 539.405 -16.835 ;
        RECT 537.715 -17.165 538.045 -16.835 ;
        RECT 536.355 -17.165 536.685 -16.835 ;
        RECT 534.995 -17.165 535.325 -16.835 ;
        RECT 533.635 -17.165 533.965 -16.835 ;
        RECT 532.275 -17.165 532.605 -16.835 ;
        RECT 530.915 -17.165 531.245 -16.835 ;
        RECT 529.555 -17.165 529.885 -16.835 ;
        RECT 528.195 -17.165 528.525 -16.835 ;
        RECT 526.835 -17.165 527.165 -16.835 ;
        RECT 525.475 -17.165 525.805 -16.835 ;
        RECT 524.115 -17.165 524.445 -16.835 ;
        RECT 522.755 -17.165 523.085 -16.835 ;
        RECT 521.395 -17.165 521.725 -16.835 ;
        RECT 520.035 -17.165 520.365 -16.835 ;
        RECT 518.675 -17.165 519.005 -16.835 ;
        RECT 517.315 -17.165 517.645 -16.835 ;
        RECT 515.955 -17.165 516.285 -16.835 ;
        RECT 514.595 -17.165 514.925 -16.835 ;
        RECT 513.235 -17.165 513.565 -16.835 ;
        RECT 511.875 -17.165 512.205 -16.835 ;
        RECT 510.515 -17.165 510.845 -16.835 ;
        RECT 509.155 -17.165 509.485 -16.835 ;
        RECT 507.795 -17.165 508.125 -16.835 ;
        RECT 506.435 -17.165 506.765 -16.835 ;
        RECT 505.075 -17.165 505.405 -16.835 ;
        RECT 503.715 -17.165 504.045 -16.835 ;
        RECT 502.355 -17.165 502.685 -16.835 ;
        RECT 500.995 -17.165 501.325 -16.835 ;
        RECT 499.635 -17.165 499.965 -16.835 ;
        RECT 498.275 -17.165 498.605 -16.835 ;
        RECT 496.915 -17.165 497.245 -16.835 ;
        RECT 495.555 -17.165 495.885 -16.835 ;
        RECT 494.195 -17.165 494.525 -16.835 ;
        RECT 492.835 -17.165 493.165 -16.835 ;
        RECT 491.475 -17.165 491.805 -16.835 ;
        RECT 490.115 -17.165 490.445 -16.835 ;
        RECT 488.755 -17.165 489.085 -16.835 ;
        RECT 487.395 -17.165 487.725 -16.835 ;
        RECT 486.035 -17.165 486.365 -16.835 ;
        RECT 484.675 -17.165 485.005 -16.835 ;
        RECT 483.315 -17.165 483.645 -16.835 ;
        RECT 481.955 -17.165 482.285 -16.835 ;
        RECT 480.595 -17.165 480.925 -16.835 ;
        RECT 479.235 -17.165 479.565 -16.835 ;
        RECT 477.875 -17.165 478.205 -16.835 ;
        RECT 476.515 -17.165 476.845 -16.835 ;
        RECT 475.155 -17.165 475.485 -16.835 ;
        RECT 473.795 -17.165 474.125 -16.835 ;
        RECT 472.435 -17.165 472.765 -16.835 ;
        RECT 471.075 -17.165 471.405 -16.835 ;
        RECT 469.715 -17.165 470.045 -16.835 ;
        RECT 468.355 -17.165 468.685 -16.835 ;
        RECT 466.995 -17.165 467.325 -16.835 ;
        RECT 465.635 -17.165 465.965 -16.835 ;
        RECT 464.275 -17.165 464.605 -16.835 ;
        RECT 462.915 -17.165 463.245 -16.835 ;
        RECT 461.555 -17.165 461.885 -16.835 ;
        RECT 460.195 -17.165 460.525 -16.835 ;
        RECT 458.835 -17.165 459.165 -16.835 ;
        RECT 457.475 -17.165 457.805 -16.835 ;
        RECT 456.115 -17.165 456.445 -16.835 ;
        RECT 454.755 -17.165 455.085 -16.835 ;
        RECT 453.395 -17.165 453.725 -16.835 ;
        RECT 452.035 -17.165 452.365 -16.835 ;
        RECT 450.675 -17.165 451.005 -16.835 ;
        RECT 449.315 -17.165 449.645 -16.835 ;
        RECT 447.955 -17.165 448.285 -16.835 ;
        RECT 446.595 -17.165 446.925 -16.835 ;
        RECT 445.235 -17.165 445.565 -16.835 ;
        RECT 443.875 -17.165 444.205 -16.835 ;
        RECT 442.515 -17.165 442.845 -16.835 ;
        RECT 441.155 -17.165 441.485 -16.835 ;
        RECT 439.795 -17.165 440.125 -16.835 ;
        RECT 438.435 -17.165 438.765 -16.835 ;
        RECT 437.075 -17.165 437.405 -16.835 ;
        RECT 435.715 -17.165 436.045 -16.835 ;
        RECT 434.355 -17.165 434.685 -16.835 ;
        RECT 432.995 -17.165 433.325 -16.835 ;
        RECT 431.635 -17.165 431.965 -16.835 ;
        RECT 430.275 -17.165 430.605 -16.835 ;
        RECT 428.915 -17.165 429.245 -16.835 ;
        RECT 427.555 -17.165 427.885 -16.835 ;
        RECT 426.195 -17.165 426.525 -16.835 ;
        RECT 424.835 -17.165 425.165 -16.835 ;
        RECT 423.475 -17.165 423.805 -16.835 ;
        RECT 422.115 -17.165 422.445 -16.835 ;
        RECT 420.755 -17.165 421.085 -16.835 ;
        RECT 419.395 -17.165 419.725 -16.835 ;
        RECT 418.035 -17.165 418.365 -16.835 ;
        RECT 416.675 -17.165 417.005 -16.835 ;
        RECT 415.315 -17.165 415.645 -16.835 ;
        RECT 413.955 -17.165 414.285 -16.835 ;
        RECT 412.595 -17.165 412.925 -16.835 ;
        RECT 411.235 -17.165 411.565 -16.835 ;
        RECT 409.875 -17.165 410.205 -16.835 ;
        RECT 408.515 -17.165 408.845 -16.835 ;
        RECT 407.155 -17.165 407.485 -16.835 ;
        RECT 405.795 -17.165 406.125 -16.835 ;
        RECT 404.435 -17.165 404.765 -16.835 ;
        RECT 403.075 -17.165 403.405 -16.835 ;
        RECT 401.715 -17.165 402.045 -16.835 ;
        RECT 400.355 -17.165 400.685 -16.835 ;
        RECT 398.995 -17.165 399.325 -16.835 ;
        RECT 397.635 -17.165 397.965 -16.835 ;
        RECT 396.275 -17.165 396.605 -16.835 ;
        RECT 394.915 -17.165 395.245 -16.835 ;
        RECT 393.555 -17.165 393.885 -16.835 ;
        RECT 392.195 -17.165 392.525 -16.835 ;
        RECT 390.835 -17.165 391.165 -16.835 ;
        RECT 389.475 -17.165 389.805 -16.835 ;
        RECT 388.115 -17.165 388.445 -16.835 ;
        RECT 386.755 -17.165 387.085 -16.835 ;
        RECT 385.395 -17.165 385.725 -16.835 ;
        RECT 384.035 -17.165 384.365 -16.835 ;
        RECT 382.675 -17.165 383.005 -16.835 ;
        RECT 381.315 -17.165 381.645 -16.835 ;
        RECT 379.955 -17.165 380.285 -16.835 ;
        RECT 378.595 -17.165 378.925 -16.835 ;
        RECT 377.235 -17.165 377.565 -16.835 ;
        RECT 375.875 -17.165 376.205 -16.835 ;
        RECT 374.515 -17.165 374.845 -16.835 ;
        RECT 373.155 -17.165 373.485 -16.835 ;
        RECT 371.795 -17.165 372.125 -16.835 ;
        RECT 370.435 -17.165 370.765 -16.835 ;
        RECT 369.075 -17.165 369.405 -16.835 ;
        RECT 367.715 -17.165 368.045 -16.835 ;
        RECT 366.355 -17.165 366.685 -16.835 ;
        RECT 364.995 -17.165 365.325 -16.835 ;
        RECT 363.635 -17.165 363.965 -16.835 ;
        RECT 362.275 -17.165 362.605 -16.835 ;
        RECT 360.915 -17.165 361.245 -16.835 ;
        RECT 359.555 -17.165 359.885 -16.835 ;
        RECT 358.195 -17.165 358.525 -16.835 ;
        RECT 356.835 -17.165 357.165 -16.835 ;
        RECT 355.475 -17.165 355.805 -16.835 ;
        RECT 354.115 -17.165 354.445 -16.835 ;
        RECT 352.755 -17.165 353.085 -16.835 ;
        RECT 351.395 -17.165 351.725 -16.835 ;
        RECT 350.035 -17.165 350.365 -16.835 ;
        RECT 348.675 -17.165 349.005 -16.835 ;
        RECT 347.315 -17.165 347.645 -16.835 ;
        RECT 345.955 -17.165 346.285 -16.835 ;
        RECT 344.595 -17.165 344.925 -16.835 ;
        RECT 343.235 -17.165 343.565 -16.835 ;
        RECT 341.875 -17.165 342.205 -16.835 ;
        RECT 340.515 -17.165 340.845 -16.835 ;
        RECT 339.155 -17.165 339.485 -16.835 ;
        RECT 337.795 -17.165 338.125 -16.835 ;
        RECT 336.435 -17.165 336.765 -16.835 ;
        RECT 335.075 -17.165 335.405 -16.835 ;
        RECT 333.715 -17.165 334.045 -16.835 ;
        RECT 332.355 -17.165 332.685 -16.835 ;
        RECT 330.995 -17.165 331.325 -16.835 ;
        RECT 329.635 -17.165 329.965 -16.835 ;
        RECT 328.275 -17.165 328.605 -16.835 ;
        RECT 326.915 -17.165 327.245 -16.835 ;
        RECT 325.555 -17.165 325.885 -16.835 ;
        RECT 324.195 -17.165 324.525 -16.835 ;
        RECT 322.835 -17.165 323.165 -16.835 ;
        RECT 321.475 -17.165 321.805 -16.835 ;
        RECT 320.115 -17.165 320.445 -16.835 ;
        RECT 318.755 -17.165 319.085 -16.835 ;
        RECT 317.395 -17.165 317.725 -16.835 ;
        RECT 316.035 -17.165 316.365 -16.835 ;
        RECT 314.675 -17.165 315.005 -16.835 ;
        RECT 313.315 -17.165 313.645 -16.835 ;
        RECT 311.955 -17.165 312.285 -16.835 ;
        RECT 310.595 -17.165 310.925 -16.835 ;
        RECT 309.235 -17.165 309.565 -16.835 ;
        RECT 307.875 -17.165 308.205 -16.835 ;
        RECT 306.515 -17.165 306.845 -16.835 ;
        RECT 305.155 -17.165 305.485 -16.835 ;
        RECT 303.795 -17.165 304.125 -16.835 ;
        RECT 302.435 -17.165 302.765 -16.835 ;
        RECT 301.075 -17.165 301.405 -16.835 ;
        RECT 299.715 -17.165 300.045 -16.835 ;
        RECT 298.355 -17.165 298.685 -16.835 ;
        RECT 296.995 -17.165 297.325 -16.835 ;
        RECT 295.635 -17.165 295.965 -16.835 ;
        RECT 294.275 -17.165 294.605 -16.835 ;
        RECT 292.915 -17.165 293.245 -16.835 ;
        RECT 291.555 -17.165 291.885 -16.835 ;
        RECT 290.195 -17.165 290.525 -16.835 ;
        RECT 288.835 -17.165 289.165 -16.835 ;
        RECT 287.475 -17.165 287.805 -16.835 ;
        RECT 286.115 -17.165 286.445 -16.835 ;
        RECT 284.755 -17.165 285.085 -16.835 ;
        RECT 283.395 -17.165 283.725 -16.835 ;
        RECT 282.035 -17.165 282.365 -16.835 ;
        RECT 280.675 -17.165 281.005 -16.835 ;
        RECT 279.315 -17.165 279.645 -16.835 ;
        RECT 277.955 -17.165 278.285 -16.835 ;
        RECT 276.595 -17.165 276.925 -16.835 ;
        RECT 275.235 -17.165 275.565 -16.835 ;
        RECT 273.875 -17.165 274.205 -16.835 ;
        RECT 272.515 -17.165 272.845 -16.835 ;
        RECT 271.155 -17.165 271.485 -16.835 ;
        RECT 269.795 -17.165 270.125 -16.835 ;
        RECT 268.435 -17.165 268.765 -16.835 ;
        RECT 267.075 -17.165 267.405 -16.835 ;
        RECT 265.715 -17.165 266.045 -16.835 ;
        RECT 264.355 -17.165 264.685 -16.835 ;
        RECT 262.995 -17.165 263.325 -16.835 ;
        RECT 261.635 -17.165 261.965 -16.835 ;
        RECT 260.275 -17.165 260.605 -16.835 ;
        RECT 258.915 -17.165 259.245 -16.835 ;
        RECT 257.555 -17.165 257.885 -16.835 ;
        RECT 256.195 -17.165 256.525 -16.835 ;
        RECT 254.835 -17.165 255.165 -16.835 ;
        RECT 253.475 -17.165 253.805 -16.835 ;
        RECT 252.115 -17.165 252.445 -16.835 ;
        RECT 250.755 -17.165 251.085 -16.835 ;
        RECT 249.395 -17.165 249.725 -16.835 ;
        RECT 248.035 -17.165 248.365 -16.835 ;
        RECT 246.675 -17.165 247.005 -16.835 ;
        RECT 245.315 -17.165 245.645 -16.835 ;
        RECT 243.955 -17.165 244.285 -16.835 ;
        RECT 242.595 -17.165 242.925 -16.835 ;
        RECT 241.235 -17.165 241.565 -16.835 ;
        RECT 239.875 -17.165 240.205 -16.835 ;
        RECT 238.515 -17.165 238.845 -16.835 ;
        RECT 237.155 -17.165 237.485 -16.835 ;
        RECT 235.795 -17.165 236.125 -16.835 ;
        RECT 234.435 -17.165 234.765 -16.835 ;
        RECT 233.075 -17.165 233.405 -16.835 ;
        RECT 231.715 -17.165 232.045 -16.835 ;
        RECT 230.355 -17.165 230.685 -16.835 ;
        RECT 228.995 -17.165 229.325 -16.835 ;
        RECT 227.635 -17.165 227.965 -16.835 ;
        RECT 226.275 -17.165 226.605 -16.835 ;
        RECT 224.915 -17.165 225.245 -16.835 ;
        RECT 223.555 -17.165 223.885 -16.835 ;
        RECT 222.195 -17.165 222.525 -16.835 ;
        RECT 220.835 -17.165 221.165 -16.835 ;
        RECT 219.475 -17.165 219.805 -16.835 ;
        RECT 218.115 -17.165 218.445 -16.835 ;
        RECT 216.755 -17.165 217.085 -16.835 ;
        RECT 215.395 -17.165 215.725 -16.835 ;
        RECT 214.035 -17.165 214.365 -16.835 ;
        RECT 212.675 -17.165 213.005 -16.835 ;
        RECT 211.315 -17.165 211.645 -16.835 ;
        RECT 209.955 -17.165 210.285 -16.835 ;
        RECT 208.595 -17.165 208.925 -16.835 ;
        RECT 207.235 -17.165 207.565 -16.835 ;
        RECT 205.875 -17.165 206.205 -16.835 ;
        RECT 204.515 -17.165 204.845 -16.835 ;
        RECT 203.155 -17.165 203.485 -16.835 ;
        RECT 201.795 -17.165 202.125 -16.835 ;
        RECT 200.435 -17.165 200.765 -16.835 ;
        RECT 199.075 -17.165 199.405 -16.835 ;
        RECT 197.715 -17.165 198.045 -16.835 ;
        RECT 196.355 -17.165 196.685 -16.835 ;
        RECT 194.995 -17.165 195.325 -16.835 ;
        RECT 193.635 -17.165 193.965 -16.835 ;
        RECT 192.275 -17.165 192.605 -16.835 ;
        RECT 190.915 -17.165 191.245 -16.835 ;
        RECT 189.555 -17.165 189.885 -16.835 ;
        RECT 188.195 -17.165 188.525 -16.835 ;
        RECT 186.835 -17.165 187.165 -16.835 ;
        RECT 185.475 -17.165 185.805 -16.835 ;
        RECT 184.115 -17.165 184.445 -16.835 ;
        RECT 182.755 -17.165 183.085 -16.835 ;
        RECT 181.395 -17.165 181.725 -16.835 ;
        RECT 180.035 -17.165 180.365 -16.835 ;
        RECT 178.675 -17.165 179.005 -16.835 ;
        RECT 177.315 -17.165 177.645 -16.835 ;
        RECT 175.955 -17.165 176.285 -16.835 ;
        RECT 174.595 -17.165 174.925 -16.835 ;
        RECT 173.235 -17.165 173.565 -16.835 ;
        RECT 171.875 -17.165 172.205 -16.835 ;
        RECT 170.515 -17.165 170.845 -16.835 ;
        RECT 169.155 -17.165 169.485 -16.835 ;
        RECT 167.795 -17.165 168.125 -16.835 ;
        RECT 166.435 -17.165 166.765 -16.835 ;
        RECT 165.075 -17.165 165.405 -16.835 ;
        RECT 163.715 -17.165 164.045 -16.835 ;
        RECT 162.355 -17.165 162.685 -16.835 ;
        RECT 160.995 -17.165 161.325 -16.835 ;
        RECT 159.635 -17.165 159.965 -16.835 ;
        RECT 158.275 -17.165 158.605 -16.835 ;
        RECT 156.915 -17.165 157.245 -16.835 ;
        RECT 155.555 -17.165 155.885 -16.835 ;
        RECT 154.195 -17.165 154.525 -16.835 ;
        RECT 152.835 -17.165 153.165 -16.835 ;
        RECT 151.475 -17.165 151.805 -16.835 ;
        RECT 150.115 -17.165 150.445 -16.835 ;
        RECT 148.755 -17.165 149.085 -16.835 ;
        RECT 147.395 -17.165 147.725 -16.835 ;
        RECT 146.035 -17.165 146.365 -16.835 ;
        RECT 144.675 -17.165 145.005 -16.835 ;
        RECT 143.315 -17.165 143.645 -16.835 ;
        RECT 141.955 -17.165 142.285 -16.835 ;
        RECT 140.595 -17.165 140.925 -16.835 ;
        RECT 139.235 -17.165 139.565 -16.835 ;
        RECT 137.875 -17.165 138.205 -16.835 ;
        RECT 136.515 -17.165 136.845 -16.835 ;
        RECT 135.155 -17.165 135.485 -16.835 ;
        RECT 133.795 -17.165 134.125 -16.835 ;
        RECT 132.435 -17.165 132.765 -16.835 ;
        RECT 131.075 -17.165 131.405 -16.835 ;
        RECT 129.715 -17.165 130.045 -16.835 ;
        RECT 128.355 -17.165 128.685 -16.835 ;
        RECT 126.995 -17.165 127.325 -16.835 ;
        RECT 125.635 -17.165 125.965 -16.835 ;
        RECT 124.275 -17.165 124.605 -16.835 ;
        RECT 678.125 -17.16 954.88 -16.84 ;
        RECT 953.875 -17.165 954.205 -16.835 ;
        RECT 952.515 -17.165 952.845 -16.835 ;
        RECT 951.155 -17.165 951.485 -16.835 ;
        RECT 949.795 -17.165 950.125 -16.835 ;
        RECT 948.435 -17.165 948.765 -16.835 ;
        RECT 947.075 -17.165 947.405 -16.835 ;
        RECT 945.715 -17.165 946.045 -16.835 ;
        RECT 944.355 -17.165 944.685 -16.835 ;
        RECT 942.995 -17.165 943.325 -16.835 ;
        RECT 941.635 -17.165 941.965 -16.835 ;
        RECT 940.275 -17.165 940.605 -16.835 ;
        RECT 938.915 -17.165 939.245 -16.835 ;
        RECT 937.555 -17.165 937.885 -16.835 ;
        RECT 936.195 -17.165 936.525 -16.835 ;
        RECT 934.835 -17.165 935.165 -16.835 ;
        RECT 933.475 -17.165 933.805 -16.835 ;
        RECT 932.115 -17.165 932.445 -16.835 ;
        RECT 930.755 -17.165 931.085 -16.835 ;
        RECT 929.395 -17.165 929.725 -16.835 ;
        RECT 928.035 -17.165 928.365 -16.835 ;
        RECT 926.675 -17.165 927.005 -16.835 ;
        RECT 925.315 -17.165 925.645 -16.835 ;
        RECT 923.955 -17.165 924.285 -16.835 ;
        RECT 922.595 -17.165 922.925 -16.835 ;
        RECT 921.235 -17.165 921.565 -16.835 ;
        RECT 919.875 -17.165 920.205 -16.835 ;
        RECT 918.515 -17.165 918.845 -16.835 ;
        RECT 917.155 -17.165 917.485 -16.835 ;
        RECT 915.795 -17.165 916.125 -16.835 ;
        RECT 914.435 -17.165 914.765 -16.835 ;
        RECT 913.075 -17.165 913.405 -16.835 ;
        RECT 911.715 -17.165 912.045 -16.835 ;
        RECT 910.355 -17.165 910.685 -16.835 ;
        RECT 908.995 -17.165 909.325 -16.835 ;
        RECT 907.635 -17.165 907.965 -16.835 ;
        RECT 906.275 -17.165 906.605 -16.835 ;
        RECT 904.915 -17.165 905.245 -16.835 ;
        RECT 903.555 -17.165 903.885 -16.835 ;
        RECT 902.195 -17.165 902.525 -16.835 ;
        RECT 900.835 -17.165 901.165 -16.835 ;
        RECT 899.475 -17.165 899.805 -16.835 ;
        RECT 898.115 -17.165 898.445 -16.835 ;
        RECT 896.755 -17.165 897.085 -16.835 ;
        RECT 895.395 -17.165 895.725 -16.835 ;
        RECT 894.035 -17.165 894.365 -16.835 ;
        RECT 892.675 -17.165 893.005 -16.835 ;
        RECT 891.315 -17.165 891.645 -16.835 ;
        RECT 889.955 -17.165 890.285 -16.835 ;
        RECT 888.595 -17.165 888.925 -16.835 ;
        RECT 887.235 -17.165 887.565 -16.835 ;
        RECT 885.875 -17.165 886.205 -16.835 ;
        RECT 884.515 -17.165 884.845 -16.835 ;
        RECT 883.155 -17.165 883.485 -16.835 ;
        RECT 881.795 -17.165 882.125 -16.835 ;
        RECT 880.435 -17.165 880.765 -16.835 ;
        RECT 879.075 -17.165 879.405 -16.835 ;
        RECT 877.715 -17.165 878.045 -16.835 ;
        RECT 876.355 -17.165 876.685 -16.835 ;
        RECT 874.995 -17.165 875.325 -16.835 ;
        RECT 873.635 -17.165 873.965 -16.835 ;
        RECT 872.275 -17.165 872.605 -16.835 ;
        RECT 870.915 -17.165 871.245 -16.835 ;
        RECT 869.555 -17.165 869.885 -16.835 ;
        RECT 868.195 -17.165 868.525 -16.835 ;
        RECT 866.835 -17.165 867.165 -16.835 ;
        RECT 865.475 -17.165 865.805 -16.835 ;
        RECT 864.115 -17.165 864.445 -16.835 ;
        RECT 862.755 -17.165 863.085 -16.835 ;
        RECT 861.395 -17.165 861.725 -16.835 ;
        RECT 860.035 -17.165 860.365 -16.835 ;
        RECT 858.675 -17.165 859.005 -16.835 ;
        RECT 857.315 -17.165 857.645 -16.835 ;
        RECT 855.955 -17.165 856.285 -16.835 ;
        RECT 854.595 -17.165 854.925 -16.835 ;
        RECT 853.235 -17.165 853.565 -16.835 ;
        RECT 851.875 -17.165 852.205 -16.835 ;
        RECT 850.515 -17.165 850.845 -16.835 ;
        RECT 849.155 -17.165 849.485 -16.835 ;
        RECT 847.795 -17.165 848.125 -16.835 ;
        RECT 846.435 -17.165 846.765 -16.835 ;
        RECT 845.075 -17.165 845.405 -16.835 ;
        RECT 843.715 -17.165 844.045 -16.835 ;
        RECT 842.355 -17.165 842.685 -16.835 ;
        RECT 840.995 -17.165 841.325 -16.835 ;
        RECT 839.635 -17.165 839.965 -16.835 ;
        RECT 838.275 -17.165 838.605 -16.835 ;
        RECT 836.915 -17.165 837.245 -16.835 ;
        RECT 835.555 -17.165 835.885 -16.835 ;
        RECT 834.195 -17.165 834.525 -16.835 ;
        RECT 832.835 -17.165 833.165 -16.835 ;
        RECT 831.475 -17.165 831.805 -16.835 ;
        RECT 830.115 -17.165 830.445 -16.835 ;
        RECT 828.755 -17.165 829.085 -16.835 ;
        RECT 827.395 -17.165 827.725 -16.835 ;
        RECT 826.035 -17.165 826.365 -16.835 ;
        RECT 824.675 -17.165 825.005 -16.835 ;
        RECT 823.315 -17.165 823.645 -16.835 ;
        RECT 821.955 -17.165 822.285 -16.835 ;
        RECT 820.595 -17.165 820.925 -16.835 ;
        RECT 819.235 -17.165 819.565 -16.835 ;
        RECT 817.875 -17.165 818.205 -16.835 ;
        RECT 816.515 -17.165 816.845 -16.835 ;
        RECT 815.155 -17.165 815.485 -16.835 ;
        RECT 813.795 -17.165 814.125 -16.835 ;
        RECT 812.435 -17.165 812.765 -16.835 ;
        RECT 811.075 -17.165 811.405 -16.835 ;
        RECT 809.715 -17.165 810.045 -16.835 ;
        RECT 808.355 -17.165 808.685 -16.835 ;
        RECT 806.995 -17.165 807.325 -16.835 ;
        RECT 805.635 -17.165 805.965 -16.835 ;
        RECT 804.275 -17.165 804.605 -16.835 ;
        RECT 802.915 -17.165 803.245 -16.835 ;
        RECT 801.555 -17.165 801.885 -16.835 ;
        RECT 800.195 -17.165 800.525 -16.835 ;
        RECT 798.835 -17.165 799.165 -16.835 ;
        RECT 797.475 -17.165 797.805 -16.835 ;
        RECT 796.115 -17.165 796.445 -16.835 ;
        RECT 794.755 -17.165 795.085 -16.835 ;
        RECT 793.395 -17.165 793.725 -16.835 ;
        RECT 792.035 -17.165 792.365 -16.835 ;
        RECT 790.675 -17.165 791.005 -16.835 ;
        RECT 789.315 -17.165 789.645 -16.835 ;
        RECT 787.955 -17.165 788.285 -16.835 ;
        RECT 786.595 -17.165 786.925 -16.835 ;
        RECT 785.235 -17.165 785.565 -16.835 ;
        RECT 783.875 -17.165 784.205 -16.835 ;
        RECT 782.515 -17.165 782.845 -16.835 ;
        RECT 781.155 -17.165 781.485 -16.835 ;
        RECT 779.795 -17.165 780.125 -16.835 ;
        RECT 778.435 -17.165 778.765 -16.835 ;
        RECT 777.075 -17.165 777.405 -16.835 ;
        RECT 775.715 -17.165 776.045 -16.835 ;
        RECT 774.355 -17.165 774.685 -16.835 ;
        RECT 772.995 -17.165 773.325 -16.835 ;
        RECT 771.635 -17.165 771.965 -16.835 ;
        RECT 770.275 -17.165 770.605 -16.835 ;
        RECT 768.915 -17.165 769.245 -16.835 ;
        RECT 767.555 -17.165 767.885 -16.835 ;
        RECT 766.195 -17.165 766.525 -16.835 ;
        RECT 764.835 -17.165 765.165 -16.835 ;
        RECT 763.475 -17.165 763.805 -16.835 ;
        RECT 762.115 -17.165 762.445 -16.835 ;
        RECT 760.755 -17.165 761.085 -16.835 ;
        RECT 759.395 -17.165 759.725 -16.835 ;
        RECT 758.035 -17.165 758.365 -16.835 ;
        RECT 756.675 -17.165 757.005 -16.835 ;
        RECT 755.315 -17.165 755.645 -16.835 ;
        RECT 753.955 -17.165 754.285 -16.835 ;
        RECT 752.595 -17.165 752.925 -16.835 ;
        RECT 751.235 -17.165 751.565 -16.835 ;
        RECT 749.875 -17.165 750.205 -16.835 ;
        RECT 748.515 -17.165 748.845 -16.835 ;
        RECT 747.155 -17.165 747.485 -16.835 ;
        RECT 745.795 -17.165 746.125 -16.835 ;
        RECT 744.435 -17.165 744.765 -16.835 ;
        RECT 743.075 -17.165 743.405 -16.835 ;
        RECT 741.715 -17.165 742.045 -16.835 ;
        RECT 740.355 -17.165 740.685 -16.835 ;
        RECT 738.995 -17.165 739.325 -16.835 ;
        RECT 737.635 -17.165 737.965 -16.835 ;
        RECT 736.275 -17.165 736.605 -16.835 ;
        RECT 734.915 -17.165 735.245 -16.835 ;
        RECT 733.555 -17.165 733.885 -16.835 ;
        RECT 732.195 -17.165 732.525 -16.835 ;
        RECT 730.835 -17.165 731.165 -16.835 ;
        RECT 729.475 -17.165 729.805 -16.835 ;
        RECT 728.115 -17.165 728.445 -16.835 ;
        RECT 726.755 -17.165 727.085 -16.835 ;
        RECT 725.395 -17.165 725.725 -16.835 ;
        RECT 724.035 -17.165 724.365 -16.835 ;
        RECT 722.675 -17.165 723.005 -16.835 ;
        RECT 721.315 -17.165 721.645 -16.835 ;
        RECT 719.955 -17.165 720.285 -16.835 ;
        RECT 718.595 -17.165 718.925 -16.835 ;
        RECT 717.235 -17.165 717.565 -16.835 ;
        RECT 715.875 -17.165 716.205 -16.835 ;
        RECT 714.515 -17.165 714.845 -16.835 ;
        RECT 713.155 -17.165 713.485 -16.835 ;
        RECT 711.795 -17.165 712.125 -16.835 ;
        RECT 710.435 -17.165 710.765 -16.835 ;
        RECT 709.075 -17.165 709.405 -16.835 ;
        RECT 707.715 -17.165 708.045 -16.835 ;
        RECT 706.355 -17.165 706.685 -16.835 ;
        RECT 704.995 -17.165 705.325 -16.835 ;
        RECT 703.635 -17.165 703.965 -16.835 ;
        RECT 702.275 -17.165 702.605 -16.835 ;
        RECT 700.915 -17.165 701.245 -16.835 ;
        RECT 699.555 -17.165 699.885 -16.835 ;
        RECT 698.195 -17.165 698.525 -16.835 ;
        RECT 696.835 -17.165 697.165 -16.835 ;
        RECT 695.475 -17.165 695.805 -16.835 ;
        RECT 694.115 -17.165 694.445 -16.835 ;
        RECT 692.755 -17.165 693.085 -16.835 ;
        RECT 691.395 -17.165 691.725 -16.835 ;
        RECT 690.035 -17.165 690.365 -16.835 ;
        RECT 688.675 -17.165 689.005 -16.835 ;
        RECT 687.315 -17.165 687.645 -16.835 ;
        RECT 685.955 -17.165 686.285 -16.835 ;
        RECT 684.595 -17.165 684.925 -16.835 ;
        RECT 683.235 -17.165 683.565 -16.835 ;
        RECT 681.875 -17.165 682.205 -16.835 ;
        RECT 680.515 -17.165 680.845 -16.835 ;
        RECT 679.155 -17.165 679.485 -16.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 -13.085 678.125 -12.755 ;
        RECT -1.52 -13.08 678.125 -12.76 ;
        RECT 676.435 -13.085 676.765 -12.755 ;
        RECT 675.075 -13.085 675.405 -12.755 ;
        RECT 673.715 -13.085 674.045 -12.755 ;
        RECT 672.355 -13.085 672.685 -12.755 ;
        RECT 670.995 -13.085 671.325 -12.755 ;
        RECT 669.635 -13.085 669.965 -12.755 ;
        RECT 668.275 -13.085 668.605 -12.755 ;
        RECT 666.915 -13.085 667.245 -12.755 ;
        RECT 665.555 -13.085 665.885 -12.755 ;
        RECT 664.195 -13.085 664.525 -12.755 ;
        RECT 662.835 -13.085 663.165 -12.755 ;
        RECT 661.475 -13.085 661.805 -12.755 ;
        RECT 660.115 -13.085 660.445 -12.755 ;
        RECT 658.755 -13.085 659.085 -12.755 ;
        RECT 657.395 -13.085 657.725 -12.755 ;
        RECT 656.035 -13.085 656.365 -12.755 ;
        RECT 654.675 -13.085 655.005 -12.755 ;
        RECT 653.315 -13.085 653.645 -12.755 ;
        RECT 651.955 -13.085 652.285 -12.755 ;
        RECT 650.595 -13.085 650.925 -12.755 ;
        RECT 649.235 -13.085 649.565 -12.755 ;
        RECT 647.875 -13.085 648.205 -12.755 ;
        RECT 646.515 -13.085 646.845 -12.755 ;
        RECT 645.155 -13.085 645.485 -12.755 ;
        RECT 643.795 -13.085 644.125 -12.755 ;
        RECT 642.435 -13.085 642.765 -12.755 ;
        RECT 641.075 -13.085 641.405 -12.755 ;
        RECT 639.715 -13.085 640.045 -12.755 ;
        RECT 638.355 -13.085 638.685 -12.755 ;
        RECT 636.995 -13.085 637.325 -12.755 ;
        RECT 635.635 -13.085 635.965 -12.755 ;
        RECT 634.275 -13.085 634.605 -12.755 ;
        RECT 632.915 -13.085 633.245 -12.755 ;
        RECT 631.555 -13.085 631.885 -12.755 ;
        RECT 630.195 -13.085 630.525 -12.755 ;
        RECT 628.835 -13.085 629.165 -12.755 ;
        RECT 627.475 -13.085 627.805 -12.755 ;
        RECT 626.115 -13.085 626.445 -12.755 ;
        RECT 624.755 -13.085 625.085 -12.755 ;
        RECT 623.395 -13.085 623.725 -12.755 ;
        RECT 622.035 -13.085 622.365 -12.755 ;
        RECT 620.675 -13.085 621.005 -12.755 ;
        RECT 619.315 -13.085 619.645 -12.755 ;
        RECT 617.955 -13.085 618.285 -12.755 ;
        RECT 616.595 -13.085 616.925 -12.755 ;
        RECT 615.235 -13.085 615.565 -12.755 ;
        RECT 613.875 -13.085 614.205 -12.755 ;
        RECT 612.515 -13.085 612.845 -12.755 ;
        RECT 611.155 -13.085 611.485 -12.755 ;
        RECT 609.795 -13.085 610.125 -12.755 ;
        RECT 608.435 -13.085 608.765 -12.755 ;
        RECT 607.075 -13.085 607.405 -12.755 ;
        RECT 605.715 -13.085 606.045 -12.755 ;
        RECT 604.355 -13.085 604.685 -12.755 ;
        RECT 602.995 -13.085 603.325 -12.755 ;
        RECT 601.635 -13.085 601.965 -12.755 ;
        RECT 600.275 -13.085 600.605 -12.755 ;
        RECT 598.915 -13.085 599.245 -12.755 ;
        RECT 597.555 -13.085 597.885 -12.755 ;
        RECT 596.195 -13.085 596.525 -12.755 ;
        RECT 594.835 -13.085 595.165 -12.755 ;
        RECT 593.475 -13.085 593.805 -12.755 ;
        RECT 592.115 -13.085 592.445 -12.755 ;
        RECT 590.755 -13.085 591.085 -12.755 ;
        RECT 589.395 -13.085 589.725 -12.755 ;
        RECT 588.035 -13.085 588.365 -12.755 ;
        RECT 586.675 -13.085 587.005 -12.755 ;
        RECT 585.315 -13.085 585.645 -12.755 ;
        RECT 583.955 -13.085 584.285 -12.755 ;
        RECT 582.595 -13.085 582.925 -12.755 ;
        RECT 581.235 -13.085 581.565 -12.755 ;
        RECT 579.875 -13.085 580.205 -12.755 ;
        RECT 578.515 -13.085 578.845 -12.755 ;
        RECT 577.155 -13.085 577.485 -12.755 ;
        RECT 575.795 -13.085 576.125 -12.755 ;
        RECT 574.435 -13.085 574.765 -12.755 ;
        RECT 573.075 -13.085 573.405 -12.755 ;
        RECT 571.715 -13.085 572.045 -12.755 ;
        RECT 570.355 -13.085 570.685 -12.755 ;
        RECT 568.995 -13.085 569.325 -12.755 ;
        RECT 567.635 -13.085 567.965 -12.755 ;
        RECT 566.275 -13.085 566.605 -12.755 ;
        RECT 564.915 -13.085 565.245 -12.755 ;
        RECT 563.555 -13.085 563.885 -12.755 ;
        RECT 562.195 -13.085 562.525 -12.755 ;
        RECT 560.835 -13.085 561.165 -12.755 ;
        RECT 559.475 -13.085 559.805 -12.755 ;
        RECT 558.115 -13.085 558.445 -12.755 ;
        RECT 556.755 -13.085 557.085 -12.755 ;
        RECT 555.395 -13.085 555.725 -12.755 ;
        RECT 554.035 -13.085 554.365 -12.755 ;
        RECT 552.675 -13.085 553.005 -12.755 ;
        RECT 551.315 -13.085 551.645 -12.755 ;
        RECT 549.955 -13.085 550.285 -12.755 ;
        RECT 548.595 -13.085 548.925 -12.755 ;
        RECT 547.235 -13.085 547.565 -12.755 ;
        RECT 545.875 -13.085 546.205 -12.755 ;
        RECT 544.515 -13.085 544.845 -12.755 ;
        RECT 543.155 -13.085 543.485 -12.755 ;
        RECT 541.795 -13.085 542.125 -12.755 ;
        RECT 540.435 -13.085 540.765 -12.755 ;
        RECT 539.075 -13.085 539.405 -12.755 ;
        RECT 537.715 -13.085 538.045 -12.755 ;
        RECT 536.355 -13.085 536.685 -12.755 ;
        RECT 534.995 -13.085 535.325 -12.755 ;
        RECT 533.635 -13.085 533.965 -12.755 ;
        RECT 532.275 -13.085 532.605 -12.755 ;
        RECT 530.915 -13.085 531.245 -12.755 ;
        RECT 529.555 -13.085 529.885 -12.755 ;
        RECT 528.195 -13.085 528.525 -12.755 ;
        RECT 526.835 -13.085 527.165 -12.755 ;
        RECT 525.475 -13.085 525.805 -12.755 ;
        RECT 524.115 -13.085 524.445 -12.755 ;
        RECT 522.755 -13.085 523.085 -12.755 ;
        RECT 521.395 -13.085 521.725 -12.755 ;
        RECT 520.035 -13.085 520.365 -12.755 ;
        RECT 518.675 -13.085 519.005 -12.755 ;
        RECT 517.315 -13.085 517.645 -12.755 ;
        RECT 515.955 -13.085 516.285 -12.755 ;
        RECT 514.595 -13.085 514.925 -12.755 ;
        RECT 513.235 -13.085 513.565 -12.755 ;
        RECT 511.875 -13.085 512.205 -12.755 ;
        RECT 510.515 -13.085 510.845 -12.755 ;
        RECT 509.155 -13.085 509.485 -12.755 ;
        RECT 507.795 -13.085 508.125 -12.755 ;
        RECT 506.435 -13.085 506.765 -12.755 ;
        RECT 505.075 -13.085 505.405 -12.755 ;
        RECT 503.715 -13.085 504.045 -12.755 ;
        RECT 502.355 -13.085 502.685 -12.755 ;
        RECT 500.995 -13.085 501.325 -12.755 ;
        RECT 499.635 -13.085 499.965 -12.755 ;
        RECT 498.275 -13.085 498.605 -12.755 ;
        RECT 496.915 -13.085 497.245 -12.755 ;
        RECT 495.555 -13.085 495.885 -12.755 ;
        RECT 494.195 -13.085 494.525 -12.755 ;
        RECT 492.835 -13.085 493.165 -12.755 ;
        RECT 491.475 -13.085 491.805 -12.755 ;
        RECT 490.115 -13.085 490.445 -12.755 ;
        RECT 488.755 -13.085 489.085 -12.755 ;
        RECT 487.395 -13.085 487.725 -12.755 ;
        RECT 486.035 -13.085 486.365 -12.755 ;
        RECT 484.675 -13.085 485.005 -12.755 ;
        RECT 483.315 -13.085 483.645 -12.755 ;
        RECT 481.955 -13.085 482.285 -12.755 ;
        RECT 480.595 -13.085 480.925 -12.755 ;
        RECT 479.235 -13.085 479.565 -12.755 ;
        RECT 477.875 -13.085 478.205 -12.755 ;
        RECT 476.515 -13.085 476.845 -12.755 ;
        RECT 475.155 -13.085 475.485 -12.755 ;
        RECT 473.795 -13.085 474.125 -12.755 ;
        RECT 472.435 -13.085 472.765 -12.755 ;
        RECT 471.075 -13.085 471.405 -12.755 ;
        RECT 469.715 -13.085 470.045 -12.755 ;
        RECT 468.355 -13.085 468.685 -12.755 ;
        RECT 466.995 -13.085 467.325 -12.755 ;
        RECT 465.635 -13.085 465.965 -12.755 ;
        RECT 464.275 -13.085 464.605 -12.755 ;
        RECT 462.915 -13.085 463.245 -12.755 ;
        RECT 461.555 -13.085 461.885 -12.755 ;
        RECT 460.195 -13.085 460.525 -12.755 ;
        RECT 458.835 -13.085 459.165 -12.755 ;
        RECT 457.475 -13.085 457.805 -12.755 ;
        RECT 456.115 -13.085 456.445 -12.755 ;
        RECT 454.755 -13.085 455.085 -12.755 ;
        RECT 453.395 -13.085 453.725 -12.755 ;
        RECT 452.035 -13.085 452.365 -12.755 ;
        RECT 450.675 -13.085 451.005 -12.755 ;
        RECT 449.315 -13.085 449.645 -12.755 ;
        RECT 447.955 -13.085 448.285 -12.755 ;
        RECT 446.595 -13.085 446.925 -12.755 ;
        RECT 445.235 -13.085 445.565 -12.755 ;
        RECT 443.875 -13.085 444.205 -12.755 ;
        RECT 442.515 -13.085 442.845 -12.755 ;
        RECT 441.155 -13.085 441.485 -12.755 ;
        RECT 439.795 -13.085 440.125 -12.755 ;
        RECT 438.435 -13.085 438.765 -12.755 ;
        RECT 437.075 -13.085 437.405 -12.755 ;
        RECT 435.715 -13.085 436.045 -12.755 ;
        RECT 434.355 -13.085 434.685 -12.755 ;
        RECT 432.995 -13.085 433.325 -12.755 ;
        RECT 431.635 -13.085 431.965 -12.755 ;
        RECT 430.275 -13.085 430.605 -12.755 ;
        RECT 428.915 -13.085 429.245 -12.755 ;
        RECT 427.555 -13.085 427.885 -12.755 ;
        RECT 426.195 -13.085 426.525 -12.755 ;
        RECT 424.835 -13.085 425.165 -12.755 ;
        RECT 423.475 -13.085 423.805 -12.755 ;
        RECT 422.115 -13.085 422.445 -12.755 ;
        RECT 420.755 -13.085 421.085 -12.755 ;
        RECT 419.395 -13.085 419.725 -12.755 ;
        RECT 418.035 -13.085 418.365 -12.755 ;
        RECT 416.675 -13.085 417.005 -12.755 ;
        RECT 415.315 -13.085 415.645 -12.755 ;
        RECT 413.955 -13.085 414.285 -12.755 ;
        RECT 412.595 -13.085 412.925 -12.755 ;
        RECT 411.235 -13.085 411.565 -12.755 ;
        RECT 409.875 -13.085 410.205 -12.755 ;
        RECT 408.515 -13.085 408.845 -12.755 ;
        RECT 407.155 -13.085 407.485 -12.755 ;
        RECT 405.795 -13.085 406.125 -12.755 ;
        RECT 404.435 -13.085 404.765 -12.755 ;
        RECT 403.075 -13.085 403.405 -12.755 ;
        RECT 401.715 -13.085 402.045 -12.755 ;
        RECT 400.355 -13.085 400.685 -12.755 ;
        RECT 398.995 -13.085 399.325 -12.755 ;
        RECT 397.635 -13.085 397.965 -12.755 ;
        RECT 396.275 -13.085 396.605 -12.755 ;
        RECT 394.915 -13.085 395.245 -12.755 ;
        RECT 393.555 -13.085 393.885 -12.755 ;
        RECT 392.195 -13.085 392.525 -12.755 ;
        RECT 390.835 -13.085 391.165 -12.755 ;
        RECT 389.475 -13.085 389.805 -12.755 ;
        RECT 388.115 -13.085 388.445 -12.755 ;
        RECT 386.755 -13.085 387.085 -12.755 ;
        RECT 385.395 -13.085 385.725 -12.755 ;
        RECT 384.035 -13.085 384.365 -12.755 ;
        RECT 382.675 -13.085 383.005 -12.755 ;
        RECT 381.315 -13.085 381.645 -12.755 ;
        RECT 379.955 -13.085 380.285 -12.755 ;
        RECT 378.595 -13.085 378.925 -12.755 ;
        RECT 377.235 -13.085 377.565 -12.755 ;
        RECT 375.875 -13.085 376.205 -12.755 ;
        RECT 374.515 -13.085 374.845 -12.755 ;
        RECT 373.155 -13.085 373.485 -12.755 ;
        RECT 371.795 -13.085 372.125 -12.755 ;
        RECT 370.435 -13.085 370.765 -12.755 ;
        RECT 369.075 -13.085 369.405 -12.755 ;
        RECT 367.715 -13.085 368.045 -12.755 ;
        RECT 366.355 -13.085 366.685 -12.755 ;
        RECT 364.995 -13.085 365.325 -12.755 ;
        RECT 363.635 -13.085 363.965 -12.755 ;
        RECT 362.275 -13.085 362.605 -12.755 ;
        RECT 360.915 -13.085 361.245 -12.755 ;
        RECT 359.555 -13.085 359.885 -12.755 ;
        RECT 358.195 -13.085 358.525 -12.755 ;
        RECT 356.835 -13.085 357.165 -12.755 ;
        RECT 355.475 -13.085 355.805 -12.755 ;
        RECT 354.115 -13.085 354.445 -12.755 ;
        RECT 352.755 -13.085 353.085 -12.755 ;
        RECT 351.395 -13.085 351.725 -12.755 ;
        RECT 350.035 -13.085 350.365 -12.755 ;
        RECT 348.675 -13.085 349.005 -12.755 ;
        RECT 347.315 -13.085 347.645 -12.755 ;
        RECT 345.955 -13.085 346.285 -12.755 ;
        RECT 344.595 -13.085 344.925 -12.755 ;
        RECT 343.235 -13.085 343.565 -12.755 ;
        RECT 341.875 -13.085 342.205 -12.755 ;
        RECT 340.515 -13.085 340.845 -12.755 ;
        RECT 339.155 -13.085 339.485 -12.755 ;
        RECT 337.795 -13.085 338.125 -12.755 ;
        RECT 336.435 -13.085 336.765 -12.755 ;
        RECT 335.075 -13.085 335.405 -12.755 ;
        RECT 333.715 -13.085 334.045 -12.755 ;
        RECT 332.355 -13.085 332.685 -12.755 ;
        RECT 330.995 -13.085 331.325 -12.755 ;
        RECT 329.635 -13.085 329.965 -12.755 ;
        RECT 328.275 -13.085 328.605 -12.755 ;
        RECT 326.915 -13.085 327.245 -12.755 ;
        RECT 325.555 -13.085 325.885 -12.755 ;
        RECT 324.195 -13.085 324.525 -12.755 ;
        RECT 322.835 -13.085 323.165 -12.755 ;
        RECT 321.475 -13.085 321.805 -12.755 ;
        RECT 320.115 -13.085 320.445 -12.755 ;
        RECT 318.755 -13.085 319.085 -12.755 ;
        RECT 317.395 -13.085 317.725 -12.755 ;
        RECT 316.035 -13.085 316.365 -12.755 ;
        RECT 314.675 -13.085 315.005 -12.755 ;
        RECT 313.315 -13.085 313.645 -12.755 ;
        RECT 311.955 -13.085 312.285 -12.755 ;
        RECT 310.595 -13.085 310.925 -12.755 ;
        RECT 309.235 -13.085 309.565 -12.755 ;
        RECT 307.875 -13.085 308.205 -12.755 ;
        RECT 306.515 -13.085 306.845 -12.755 ;
        RECT 305.155 -13.085 305.485 -12.755 ;
        RECT 303.795 -13.085 304.125 -12.755 ;
        RECT 302.435 -13.085 302.765 -12.755 ;
        RECT 301.075 -13.085 301.405 -12.755 ;
        RECT 299.715 -13.085 300.045 -12.755 ;
        RECT 298.355 -13.085 298.685 -12.755 ;
        RECT 296.995 -13.085 297.325 -12.755 ;
        RECT 295.635 -13.085 295.965 -12.755 ;
        RECT 294.275 -13.085 294.605 -12.755 ;
        RECT 292.915 -13.085 293.245 -12.755 ;
        RECT 291.555 -13.085 291.885 -12.755 ;
        RECT 290.195 -13.085 290.525 -12.755 ;
        RECT 288.835 -13.085 289.165 -12.755 ;
        RECT 287.475 -13.085 287.805 -12.755 ;
        RECT 286.115 -13.085 286.445 -12.755 ;
        RECT 284.755 -13.085 285.085 -12.755 ;
        RECT 283.395 -13.085 283.725 -12.755 ;
        RECT 282.035 -13.085 282.365 -12.755 ;
        RECT 280.675 -13.085 281.005 -12.755 ;
        RECT 279.315 -13.085 279.645 -12.755 ;
        RECT 277.955 -13.085 278.285 -12.755 ;
        RECT 276.595 -13.085 276.925 -12.755 ;
        RECT 275.235 -13.085 275.565 -12.755 ;
        RECT 273.875 -13.085 274.205 -12.755 ;
        RECT 272.515 -13.085 272.845 -12.755 ;
        RECT 271.155 -13.085 271.485 -12.755 ;
        RECT 269.795 -13.085 270.125 -12.755 ;
        RECT 268.435 -13.085 268.765 -12.755 ;
        RECT 267.075 -13.085 267.405 -12.755 ;
        RECT 265.715 -13.085 266.045 -12.755 ;
        RECT 264.355 -13.085 264.685 -12.755 ;
        RECT 262.995 -13.085 263.325 -12.755 ;
        RECT 261.635 -13.085 261.965 -12.755 ;
        RECT 260.275 -13.085 260.605 -12.755 ;
        RECT 258.915 -13.085 259.245 -12.755 ;
        RECT 257.555 -13.085 257.885 -12.755 ;
        RECT 256.195 -13.085 256.525 -12.755 ;
        RECT 254.835 -13.085 255.165 -12.755 ;
        RECT 253.475 -13.085 253.805 -12.755 ;
        RECT 252.115 -13.085 252.445 -12.755 ;
        RECT 250.755 -13.085 251.085 -12.755 ;
        RECT 249.395 -13.085 249.725 -12.755 ;
        RECT 248.035 -13.085 248.365 -12.755 ;
        RECT 246.675 -13.085 247.005 -12.755 ;
        RECT 245.315 -13.085 245.645 -12.755 ;
        RECT 243.955 -13.085 244.285 -12.755 ;
        RECT 242.595 -13.085 242.925 -12.755 ;
        RECT 241.235 -13.085 241.565 -12.755 ;
        RECT 239.875 -13.085 240.205 -12.755 ;
        RECT 238.515 -13.085 238.845 -12.755 ;
        RECT 237.155 -13.085 237.485 -12.755 ;
        RECT 235.795 -13.085 236.125 -12.755 ;
        RECT 234.435 -13.085 234.765 -12.755 ;
        RECT 233.075 -13.085 233.405 -12.755 ;
        RECT 231.715 -13.085 232.045 -12.755 ;
        RECT 230.355 -13.085 230.685 -12.755 ;
        RECT 228.995 -13.085 229.325 -12.755 ;
        RECT 227.635 -13.085 227.965 -12.755 ;
        RECT 226.275 -13.085 226.605 -12.755 ;
        RECT 224.915 -13.085 225.245 -12.755 ;
        RECT 223.555 -13.085 223.885 -12.755 ;
        RECT 222.195 -13.085 222.525 -12.755 ;
        RECT 220.835 -13.085 221.165 -12.755 ;
        RECT 219.475 -13.085 219.805 -12.755 ;
        RECT 218.115 -13.085 218.445 -12.755 ;
        RECT 216.755 -13.085 217.085 -12.755 ;
        RECT 215.395 -13.085 215.725 -12.755 ;
        RECT 214.035 -13.085 214.365 -12.755 ;
        RECT 212.675 -13.085 213.005 -12.755 ;
        RECT 211.315 -13.085 211.645 -12.755 ;
        RECT 209.955 -13.085 210.285 -12.755 ;
        RECT 208.595 -13.085 208.925 -12.755 ;
        RECT 207.235 -13.085 207.565 -12.755 ;
        RECT 205.875 -13.085 206.205 -12.755 ;
        RECT 204.515 -13.085 204.845 -12.755 ;
        RECT 203.155 -13.085 203.485 -12.755 ;
        RECT 201.795 -13.085 202.125 -12.755 ;
        RECT 200.435 -13.085 200.765 -12.755 ;
        RECT 199.075 -13.085 199.405 -12.755 ;
        RECT 197.715 -13.085 198.045 -12.755 ;
        RECT 196.355 -13.085 196.685 -12.755 ;
        RECT 194.995 -13.085 195.325 -12.755 ;
        RECT 193.635 -13.085 193.965 -12.755 ;
        RECT 192.275 -13.085 192.605 -12.755 ;
        RECT 190.915 -13.085 191.245 -12.755 ;
        RECT 189.555 -13.085 189.885 -12.755 ;
        RECT 188.195 -13.085 188.525 -12.755 ;
        RECT 186.835 -13.085 187.165 -12.755 ;
        RECT 185.475 -13.085 185.805 -12.755 ;
        RECT 184.115 -13.085 184.445 -12.755 ;
        RECT 182.755 -13.085 183.085 -12.755 ;
        RECT 181.395 -13.085 181.725 -12.755 ;
        RECT 180.035 -13.085 180.365 -12.755 ;
        RECT 178.675 -13.085 179.005 -12.755 ;
        RECT 177.315 -13.085 177.645 -12.755 ;
        RECT 175.955 -13.085 176.285 -12.755 ;
        RECT 174.595 -13.085 174.925 -12.755 ;
        RECT 173.235 -13.085 173.565 -12.755 ;
        RECT 171.875 -13.085 172.205 -12.755 ;
        RECT 170.515 -13.085 170.845 -12.755 ;
        RECT 169.155 -13.085 169.485 -12.755 ;
        RECT 167.795 -13.085 168.125 -12.755 ;
        RECT 166.435 -13.085 166.765 -12.755 ;
        RECT 165.075 -13.085 165.405 -12.755 ;
        RECT 163.715 -13.085 164.045 -12.755 ;
        RECT 162.355 -13.085 162.685 -12.755 ;
        RECT 160.995 -13.085 161.325 -12.755 ;
        RECT 159.635 -13.085 159.965 -12.755 ;
        RECT 158.275 -13.085 158.605 -12.755 ;
        RECT 156.915 -13.085 157.245 -12.755 ;
        RECT 155.555 -13.085 155.885 -12.755 ;
        RECT 154.195 -13.085 154.525 -12.755 ;
        RECT 152.835 -13.085 153.165 -12.755 ;
        RECT 151.475 -13.085 151.805 -12.755 ;
        RECT 150.115 -13.085 150.445 -12.755 ;
        RECT 148.755 -13.085 149.085 -12.755 ;
        RECT 147.395 -13.085 147.725 -12.755 ;
        RECT 146.035 -13.085 146.365 -12.755 ;
        RECT 144.675 -13.085 145.005 -12.755 ;
        RECT 143.315 -13.085 143.645 -12.755 ;
        RECT 141.955 -13.085 142.285 -12.755 ;
        RECT 140.595 -13.085 140.925 -12.755 ;
        RECT 139.235 -13.085 139.565 -12.755 ;
        RECT 137.875 -13.085 138.205 -12.755 ;
        RECT 136.515 -13.085 136.845 -12.755 ;
        RECT 135.155 -13.085 135.485 -12.755 ;
        RECT 133.795 -13.085 134.125 -12.755 ;
        RECT 132.435 -13.085 132.765 -12.755 ;
        RECT 131.075 -13.085 131.405 -12.755 ;
        RECT 129.715 -13.085 130.045 -12.755 ;
        RECT 128.355 -13.085 128.685 -12.755 ;
        RECT 126.995 -13.085 127.325 -12.755 ;
        RECT 125.635 -13.085 125.965 -12.755 ;
        RECT 124.275 -13.085 124.605 -12.755 ;
        RECT 122.915 -13.085 123.245 -12.755 ;
        RECT 121.555 -13.085 121.885 -12.755 ;
        RECT 120.195 -13.085 120.525 -12.755 ;
        RECT 118.835 -13.085 119.165 -12.755 ;
        RECT 117.475 -13.085 117.805 -12.755 ;
        RECT 116.115 -13.085 116.445 -12.755 ;
        RECT 114.755 -13.085 115.085 -12.755 ;
        RECT 113.395 -13.085 113.725 -12.755 ;
        RECT 112.035 -13.085 112.365 -12.755 ;
        RECT 110.675 -13.085 111.005 -12.755 ;
        RECT 109.315 -13.085 109.645 -12.755 ;
        RECT 107.955 -13.085 108.285 -12.755 ;
        RECT 106.595 -13.085 106.925 -12.755 ;
        RECT 105.235 -13.085 105.565 -12.755 ;
        RECT 103.875 -13.085 104.205 -12.755 ;
        RECT 102.515 -13.085 102.845 -12.755 ;
        RECT 101.155 -13.085 101.485 -12.755 ;
        RECT 99.795 -13.085 100.125 -12.755 ;
        RECT 98.435 -13.085 98.765 -12.755 ;
        RECT 97.075 -13.085 97.405 -12.755 ;
        RECT 95.715 -13.085 96.045 -12.755 ;
        RECT 94.355 -13.085 94.685 -12.755 ;
        RECT 92.995 -13.085 93.325 -12.755 ;
        RECT 91.635 -13.085 91.965 -12.755 ;
        RECT 90.275 -13.085 90.605 -12.755 ;
        RECT 88.915 -13.085 89.245 -12.755 ;
        RECT 87.555 -13.085 87.885 -12.755 ;
        RECT 86.195 -13.085 86.525 -12.755 ;
        RECT 84.835 -13.085 85.165 -12.755 ;
        RECT 83.475 -13.085 83.805 -12.755 ;
        RECT 82.115 -13.085 82.445 -12.755 ;
        RECT 80.755 -13.085 81.085 -12.755 ;
        RECT 79.395 -13.085 79.725 -12.755 ;
        RECT 78.035 -13.085 78.365 -12.755 ;
        RECT 76.675 -13.085 77.005 -12.755 ;
        RECT 75.315 -13.085 75.645 -12.755 ;
        RECT 73.955 -13.085 74.285 -12.755 ;
        RECT 72.595 -13.085 72.925 -12.755 ;
        RECT 71.235 -13.085 71.565 -12.755 ;
        RECT 69.875 -13.085 70.205 -12.755 ;
        RECT 68.515 -13.085 68.845 -12.755 ;
        RECT 67.155 -13.085 67.485 -12.755 ;
        RECT 65.795 -13.085 66.125 -12.755 ;
        RECT 64.435 -13.085 64.765 -12.755 ;
        RECT 63.075 -13.085 63.405 -12.755 ;
        RECT 61.715 -13.085 62.045 -12.755 ;
        RECT 60.355 -13.085 60.685 -12.755 ;
        RECT 58.995 -13.085 59.325 -12.755 ;
        RECT 57.635 -13.085 57.965 -12.755 ;
        RECT 56.275 -13.085 56.605 -12.755 ;
        RECT 54.915 -13.085 55.245 -12.755 ;
        RECT 53.555 -13.085 53.885 -12.755 ;
        RECT 52.195 -13.085 52.525 -12.755 ;
        RECT 50.835 -13.085 51.165 -12.755 ;
        RECT 49.475 -13.085 49.805 -12.755 ;
        RECT 48.115 -13.085 48.445 -12.755 ;
        RECT 46.755 -13.085 47.085 -12.755 ;
        RECT 45.395 -13.085 45.725 -12.755 ;
        RECT 44.035 -13.085 44.365 -12.755 ;
        RECT 42.675 -13.085 43.005 -12.755 ;
        RECT 41.315 -13.085 41.645 -12.755 ;
        RECT 39.955 -13.085 40.285 -12.755 ;
        RECT 38.595 -13.085 38.925 -12.755 ;
        RECT 37.235 -13.085 37.565 -12.755 ;
        RECT 35.875 -13.085 36.205 -12.755 ;
        RECT 34.515 -13.085 34.845 -12.755 ;
        RECT 33.155 -13.085 33.485 -12.755 ;
        RECT 31.795 -13.085 32.125 -12.755 ;
        RECT 30.435 -13.085 30.765 -12.755 ;
        RECT 29.075 -13.085 29.405 -12.755 ;
        RECT 27.715 -13.085 28.045 -12.755 ;
        RECT 26.355 -13.085 26.685 -12.755 ;
        RECT 24.995 -13.085 25.325 -12.755 ;
        RECT 23.635 -13.085 23.965 -12.755 ;
        RECT 22.275 -13.085 22.605 -12.755 ;
        RECT 20.915 -13.085 21.245 -12.755 ;
        RECT 19.555 -13.085 19.885 -12.755 ;
        RECT 18.195 -13.085 18.525 -12.755 ;
        RECT 16.835 -13.085 17.165 -12.755 ;
        RECT 15.475 -13.085 15.805 -12.755 ;
        RECT 14.115 -13.085 14.445 -12.755 ;
        RECT 12.755 -13.085 13.085 -12.755 ;
        RECT 11.395 -13.085 11.725 -12.755 ;
        RECT 10.035 -13.085 10.365 -12.755 ;
        RECT 8.675 -13.085 9.005 -12.755 ;
        RECT 7.315 -13.085 7.645 -12.755 ;
        RECT 5.955 -13.085 6.285 -12.755 ;
        RECT 4.595 -13.085 4.925 -12.755 ;
        RECT 3.235 -13.085 3.565 -12.755 ;
        RECT 1.875 -13.085 2.205 -12.755 ;
        RECT 0.515 -13.085 0.845 -12.755 ;
        RECT -0.845 -13.085 -0.515 -12.755 ;
        RECT 678.125 -13.08 954.88 -12.76 ;
        RECT 953.875 -13.085 954.205 -12.755 ;
        RECT 952.515 -13.085 952.845 -12.755 ;
        RECT 951.155 -13.085 951.485 -12.755 ;
        RECT 949.795 -13.085 950.125 -12.755 ;
        RECT 948.435 -13.085 948.765 -12.755 ;
        RECT 947.075 -13.085 947.405 -12.755 ;
        RECT 945.715 -13.085 946.045 -12.755 ;
        RECT 944.355 -13.085 944.685 -12.755 ;
        RECT 942.995 -13.085 943.325 -12.755 ;
        RECT 941.635 -13.085 941.965 -12.755 ;
        RECT 940.275 -13.085 940.605 -12.755 ;
        RECT 938.915 -13.085 939.245 -12.755 ;
        RECT 937.555 -13.085 937.885 -12.755 ;
        RECT 936.195 -13.085 936.525 -12.755 ;
        RECT 934.835 -13.085 935.165 -12.755 ;
        RECT 933.475 -13.085 933.805 -12.755 ;
        RECT 932.115 -13.085 932.445 -12.755 ;
        RECT 930.755 -13.085 931.085 -12.755 ;
        RECT 929.395 -13.085 929.725 -12.755 ;
        RECT 928.035 -13.085 928.365 -12.755 ;
        RECT 926.675 -13.085 927.005 -12.755 ;
        RECT 925.315 -13.085 925.645 -12.755 ;
        RECT 923.955 -13.085 924.285 -12.755 ;
        RECT 922.595 -13.085 922.925 -12.755 ;
        RECT 921.235 -13.085 921.565 -12.755 ;
        RECT 919.875 -13.085 920.205 -12.755 ;
        RECT 918.515 -13.085 918.845 -12.755 ;
        RECT 917.155 -13.085 917.485 -12.755 ;
        RECT 915.795 -13.085 916.125 -12.755 ;
        RECT 914.435 -13.085 914.765 -12.755 ;
        RECT 913.075 -13.085 913.405 -12.755 ;
        RECT 911.715 -13.085 912.045 -12.755 ;
        RECT 910.355 -13.085 910.685 -12.755 ;
        RECT 908.995 -13.085 909.325 -12.755 ;
        RECT 907.635 -13.085 907.965 -12.755 ;
        RECT 906.275 -13.085 906.605 -12.755 ;
        RECT 904.915 -13.085 905.245 -12.755 ;
        RECT 903.555 -13.085 903.885 -12.755 ;
        RECT 902.195 -13.085 902.525 -12.755 ;
        RECT 900.835 -13.085 901.165 -12.755 ;
        RECT 899.475 -13.085 899.805 -12.755 ;
        RECT 898.115 -13.085 898.445 -12.755 ;
        RECT 896.755 -13.085 897.085 -12.755 ;
        RECT 895.395 -13.085 895.725 -12.755 ;
        RECT 894.035 -13.085 894.365 -12.755 ;
        RECT 892.675 -13.085 893.005 -12.755 ;
        RECT 891.315 -13.085 891.645 -12.755 ;
        RECT 889.955 -13.085 890.285 -12.755 ;
        RECT 888.595 -13.085 888.925 -12.755 ;
        RECT 887.235 -13.085 887.565 -12.755 ;
        RECT 885.875 -13.085 886.205 -12.755 ;
        RECT 884.515 -13.085 884.845 -12.755 ;
        RECT 883.155 -13.085 883.485 -12.755 ;
        RECT 881.795 -13.085 882.125 -12.755 ;
        RECT 880.435 -13.085 880.765 -12.755 ;
        RECT 879.075 -13.085 879.405 -12.755 ;
        RECT 877.715 -13.085 878.045 -12.755 ;
        RECT 876.355 -13.085 876.685 -12.755 ;
        RECT 874.995 -13.085 875.325 -12.755 ;
        RECT 873.635 -13.085 873.965 -12.755 ;
        RECT 872.275 -13.085 872.605 -12.755 ;
        RECT 870.915 -13.085 871.245 -12.755 ;
        RECT 869.555 -13.085 869.885 -12.755 ;
        RECT 868.195 -13.085 868.525 -12.755 ;
        RECT 866.835 -13.085 867.165 -12.755 ;
        RECT 865.475 -13.085 865.805 -12.755 ;
        RECT 864.115 -13.085 864.445 -12.755 ;
        RECT 862.755 -13.085 863.085 -12.755 ;
        RECT 861.395 -13.085 861.725 -12.755 ;
        RECT 860.035 -13.085 860.365 -12.755 ;
        RECT 858.675 -13.085 859.005 -12.755 ;
        RECT 857.315 -13.085 857.645 -12.755 ;
        RECT 855.955 -13.085 856.285 -12.755 ;
        RECT 854.595 -13.085 854.925 -12.755 ;
        RECT 853.235 -13.085 853.565 -12.755 ;
        RECT 851.875 -13.085 852.205 -12.755 ;
        RECT 850.515 -13.085 850.845 -12.755 ;
        RECT 849.155 -13.085 849.485 -12.755 ;
        RECT 847.795 -13.085 848.125 -12.755 ;
        RECT 846.435 -13.085 846.765 -12.755 ;
        RECT 845.075 -13.085 845.405 -12.755 ;
        RECT 843.715 -13.085 844.045 -12.755 ;
        RECT 842.355 -13.085 842.685 -12.755 ;
        RECT 840.995 -13.085 841.325 -12.755 ;
        RECT 839.635 -13.085 839.965 -12.755 ;
        RECT 838.275 -13.085 838.605 -12.755 ;
        RECT 836.915 -13.085 837.245 -12.755 ;
        RECT 835.555 -13.085 835.885 -12.755 ;
        RECT 834.195 -13.085 834.525 -12.755 ;
        RECT 832.835 -13.085 833.165 -12.755 ;
        RECT 831.475 -13.085 831.805 -12.755 ;
        RECT 830.115 -13.085 830.445 -12.755 ;
        RECT 828.755 -13.085 829.085 -12.755 ;
        RECT 827.395 -13.085 827.725 -12.755 ;
        RECT 826.035 -13.085 826.365 -12.755 ;
        RECT 824.675 -13.085 825.005 -12.755 ;
        RECT 823.315 -13.085 823.645 -12.755 ;
        RECT 821.955 -13.085 822.285 -12.755 ;
        RECT 820.595 -13.085 820.925 -12.755 ;
        RECT 819.235 -13.085 819.565 -12.755 ;
        RECT 817.875 -13.085 818.205 -12.755 ;
        RECT 816.515 -13.085 816.845 -12.755 ;
        RECT 815.155 -13.085 815.485 -12.755 ;
        RECT 813.795 -13.085 814.125 -12.755 ;
        RECT 812.435 -13.085 812.765 -12.755 ;
        RECT 811.075 -13.085 811.405 -12.755 ;
        RECT 809.715 -13.085 810.045 -12.755 ;
        RECT 808.355 -13.085 808.685 -12.755 ;
        RECT 806.995 -13.085 807.325 -12.755 ;
        RECT 805.635 -13.085 805.965 -12.755 ;
        RECT 804.275 -13.085 804.605 -12.755 ;
        RECT 802.915 -13.085 803.245 -12.755 ;
        RECT 801.555 -13.085 801.885 -12.755 ;
        RECT 800.195 -13.085 800.525 -12.755 ;
        RECT 798.835 -13.085 799.165 -12.755 ;
        RECT 797.475 -13.085 797.805 -12.755 ;
        RECT 796.115 -13.085 796.445 -12.755 ;
        RECT 794.755 -13.085 795.085 -12.755 ;
        RECT 793.395 -13.085 793.725 -12.755 ;
        RECT 792.035 -13.085 792.365 -12.755 ;
        RECT 790.675 -13.085 791.005 -12.755 ;
        RECT 789.315 -13.085 789.645 -12.755 ;
        RECT 787.955 -13.085 788.285 -12.755 ;
        RECT 786.595 -13.085 786.925 -12.755 ;
        RECT 785.235 -13.085 785.565 -12.755 ;
        RECT 783.875 -13.085 784.205 -12.755 ;
        RECT 782.515 -13.085 782.845 -12.755 ;
        RECT 781.155 -13.085 781.485 -12.755 ;
        RECT 779.795 -13.085 780.125 -12.755 ;
        RECT 778.435 -13.085 778.765 -12.755 ;
        RECT 777.075 -13.085 777.405 -12.755 ;
        RECT 775.715 -13.085 776.045 -12.755 ;
        RECT 774.355 -13.085 774.685 -12.755 ;
        RECT 772.995 -13.085 773.325 -12.755 ;
        RECT 771.635 -13.085 771.965 -12.755 ;
        RECT 770.275 -13.085 770.605 -12.755 ;
        RECT 768.915 -13.085 769.245 -12.755 ;
        RECT 767.555 -13.085 767.885 -12.755 ;
        RECT 766.195 -13.085 766.525 -12.755 ;
        RECT 764.835 -13.085 765.165 -12.755 ;
        RECT 763.475 -13.085 763.805 -12.755 ;
        RECT 762.115 -13.085 762.445 -12.755 ;
        RECT 760.755 -13.085 761.085 -12.755 ;
        RECT 759.395 -13.085 759.725 -12.755 ;
        RECT 758.035 -13.085 758.365 -12.755 ;
        RECT 756.675 -13.085 757.005 -12.755 ;
        RECT 755.315 -13.085 755.645 -12.755 ;
        RECT 753.955 -13.085 754.285 -12.755 ;
        RECT 752.595 -13.085 752.925 -12.755 ;
        RECT 751.235 -13.085 751.565 -12.755 ;
        RECT 749.875 -13.085 750.205 -12.755 ;
        RECT 748.515 -13.085 748.845 -12.755 ;
        RECT 747.155 -13.085 747.485 -12.755 ;
        RECT 745.795 -13.085 746.125 -12.755 ;
        RECT 744.435 -13.085 744.765 -12.755 ;
        RECT 743.075 -13.085 743.405 -12.755 ;
        RECT 741.715 -13.085 742.045 -12.755 ;
        RECT 740.355 -13.085 740.685 -12.755 ;
        RECT 738.995 -13.085 739.325 -12.755 ;
        RECT 737.635 -13.085 737.965 -12.755 ;
        RECT 736.275 -13.085 736.605 -12.755 ;
        RECT 734.915 -13.085 735.245 -12.755 ;
        RECT 733.555 -13.085 733.885 -12.755 ;
        RECT 732.195 -13.085 732.525 -12.755 ;
        RECT 730.835 -13.085 731.165 -12.755 ;
        RECT 729.475 -13.085 729.805 -12.755 ;
        RECT 728.115 -13.085 728.445 -12.755 ;
        RECT 726.755 -13.085 727.085 -12.755 ;
        RECT 725.395 -13.085 725.725 -12.755 ;
        RECT 724.035 -13.085 724.365 -12.755 ;
        RECT 722.675 -13.085 723.005 -12.755 ;
        RECT 721.315 -13.085 721.645 -12.755 ;
        RECT 719.955 -13.085 720.285 -12.755 ;
        RECT 718.595 -13.085 718.925 -12.755 ;
        RECT 717.235 -13.085 717.565 -12.755 ;
        RECT 715.875 -13.085 716.205 -12.755 ;
        RECT 714.515 -13.085 714.845 -12.755 ;
        RECT 713.155 -13.085 713.485 -12.755 ;
        RECT 711.795 -13.085 712.125 -12.755 ;
        RECT 710.435 -13.085 710.765 -12.755 ;
        RECT 709.075 -13.085 709.405 -12.755 ;
        RECT 707.715 -13.085 708.045 -12.755 ;
        RECT 706.355 -13.085 706.685 -12.755 ;
        RECT 704.995 -13.085 705.325 -12.755 ;
        RECT 703.635 -13.085 703.965 -12.755 ;
        RECT 702.275 -13.085 702.605 -12.755 ;
        RECT 700.915 -13.085 701.245 -12.755 ;
        RECT 699.555 -13.085 699.885 -12.755 ;
        RECT 698.195 -13.085 698.525 -12.755 ;
        RECT 696.835 -13.085 697.165 -12.755 ;
        RECT 695.475 -13.085 695.805 -12.755 ;
        RECT 694.115 -13.085 694.445 -12.755 ;
        RECT 692.755 -13.085 693.085 -12.755 ;
        RECT 691.395 -13.085 691.725 -12.755 ;
        RECT 690.035 -13.085 690.365 -12.755 ;
        RECT 688.675 -13.085 689.005 -12.755 ;
        RECT 687.315 -13.085 687.645 -12.755 ;
        RECT 685.955 -13.085 686.285 -12.755 ;
        RECT 684.595 -13.085 684.925 -12.755 ;
        RECT 683.235 -13.085 683.565 -12.755 ;
        RECT 681.875 -13.085 682.205 -12.755 ;
        RECT 680.515 -13.085 680.845 -12.755 ;
        RECT 679.155 -13.085 679.485 -12.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 -14.445 125.965 -14.115 ;
        RECT 124.275 -14.445 124.605 -14.115 ;
        RECT 122.915 -14.445 123.245 -14.115 ;
        RECT 121.555 -14.445 121.885 -14.115 ;
        RECT 120.195 -14.445 120.525 -14.115 ;
        RECT 118.835 -14.445 119.165 -14.115 ;
        RECT 117.475 -14.445 117.805 -14.115 ;
        RECT 116.115 -14.445 116.445 -14.115 ;
        RECT 114.755 -14.445 115.085 -14.115 ;
        RECT 113.395 -14.445 113.725 -14.115 ;
        RECT 112.035 -14.445 112.365 -14.115 ;
        RECT 110.675 -14.445 111.005 -14.115 ;
        RECT 109.315 -14.445 109.645 -14.115 ;
        RECT 107.955 -14.445 108.285 -14.115 ;
        RECT 106.595 -14.445 106.925 -14.115 ;
        RECT 105.235 -14.445 105.565 -14.115 ;
        RECT 103.875 -14.445 104.205 -14.115 ;
        RECT 102.515 -14.445 102.845 -14.115 ;
        RECT 101.155 -14.445 101.485 -14.115 ;
        RECT 99.795 -14.445 100.125 -14.115 ;
        RECT 98.435 -14.445 98.765 -14.115 ;
        RECT 97.075 -14.445 97.405 -14.115 ;
        RECT 95.715 -14.445 96.045 -14.115 ;
        RECT 94.355 -14.445 94.685 -14.115 ;
        RECT 92.995 -14.445 93.325 -14.115 ;
        RECT 91.635 -14.445 91.965 -14.115 ;
        RECT 90.275 -14.445 90.605 -14.115 ;
        RECT 88.915 -14.445 89.245 -14.115 ;
        RECT 87.555 -14.445 87.885 -14.115 ;
        RECT 86.195 -14.445 86.525 -14.115 ;
        RECT 84.835 -14.445 85.165 -14.115 ;
        RECT 83.475 -14.445 83.805 -14.115 ;
        RECT 82.115 -14.445 82.445 -14.115 ;
        RECT 80.755 -14.445 81.085 -14.115 ;
        RECT 79.395 -14.445 79.725 -14.115 ;
        RECT 78.035 -14.445 78.365 -14.115 ;
        RECT 76.675 -14.445 77.005 -14.115 ;
        RECT 75.315 -14.445 75.645 -14.115 ;
        RECT 73.955 -14.445 74.285 -14.115 ;
        RECT 72.595 -14.445 72.925 -14.115 ;
        RECT 71.235 -14.445 71.565 -14.115 ;
        RECT 69.875 -14.445 70.205 -14.115 ;
        RECT 68.515 -14.445 68.845 -14.115 ;
        RECT 67.155 -14.445 67.485 -14.115 ;
        RECT 65.795 -14.445 66.125 -14.115 ;
        RECT 64.435 -14.445 64.765 -14.115 ;
        RECT 63.075 -14.445 63.405 -14.115 ;
        RECT 61.715 -14.445 62.045 -14.115 ;
        RECT 60.355 -14.445 60.685 -14.115 ;
        RECT 58.995 -14.445 59.325 -14.115 ;
        RECT 57.635 -14.445 57.965 -14.115 ;
        RECT 56.275 -14.445 56.605 -14.115 ;
        RECT 54.915 -14.445 55.245 -14.115 ;
        RECT 53.555 -14.445 53.885 -14.115 ;
        RECT 52.195 -14.445 52.525 -14.115 ;
        RECT 50.835 -14.445 51.165 -14.115 ;
        RECT 49.475 -14.445 49.805 -14.115 ;
        RECT 48.115 -14.445 48.445 -14.115 ;
        RECT 46.755 -14.445 47.085 -14.115 ;
        RECT 45.395 -14.445 45.725 -14.115 ;
        RECT 44.035 -14.445 44.365 -14.115 ;
        RECT 42.675 -14.445 43.005 -14.115 ;
        RECT 41.315 -14.445 41.645 -14.115 ;
        RECT 39.955 -14.445 40.285 -14.115 ;
        RECT 38.595 -14.445 38.925 -14.115 ;
        RECT 37.235 -14.445 37.565 -14.115 ;
        RECT 35.875 -14.445 36.205 -14.115 ;
        RECT 34.515 -14.445 34.845 -14.115 ;
        RECT 33.155 -14.445 33.485 -14.115 ;
        RECT 31.795 -14.445 32.125 -14.115 ;
        RECT 30.435 -14.445 30.765 -14.115 ;
        RECT 29.075 -14.445 29.405 -14.115 ;
        RECT 27.715 -14.445 28.045 -14.115 ;
        RECT 26.355 -14.445 26.685 -14.115 ;
        RECT 24.995 -14.445 25.325 -14.115 ;
        RECT 23.635 -14.445 23.965 -14.115 ;
        RECT 22.275 -14.445 22.605 -14.115 ;
        RECT 20.915 -14.445 21.245 -14.115 ;
        RECT 19.555 -14.445 19.885 -14.115 ;
        RECT 18.195 -14.445 18.525 -14.115 ;
        RECT 16.835 -14.445 17.165 -14.115 ;
        RECT 15.475 -14.445 15.805 -14.115 ;
        RECT 14.115 -14.445 14.445 -14.115 ;
        RECT 12.755 -14.445 13.085 -14.115 ;
        RECT 11.395 -14.445 11.725 -14.115 ;
        RECT 10.035 -14.445 10.365 -14.115 ;
        RECT 8.675 -14.445 9.005 -14.115 ;
        RECT 7.315 -14.445 7.645 -14.115 ;
        RECT 5.955 -14.445 6.285 -14.115 ;
        RECT 4.595 -14.445 4.925 -14.115 ;
        RECT 3.235 -14.445 3.565 -14.115 ;
        RECT 1.875 -14.445 2.205 -14.115 ;
        RECT 0.515 -14.445 0.845 -14.115 ;
        RECT -0.845 -14.445 -0.515 -14.115 ;
        RECT 677.795 -14.445 678.125 -14.115 ;
        RECT -1.52 -14.44 678.125 -14.12 ;
        RECT 676.435 -14.445 676.765 -14.115 ;
        RECT 675.075 -14.445 675.405 -14.115 ;
        RECT 673.715 -14.445 674.045 -14.115 ;
        RECT 672.355 -14.445 672.685 -14.115 ;
        RECT 670.995 -14.445 671.325 -14.115 ;
        RECT 669.635 -14.445 669.965 -14.115 ;
        RECT 668.275 -14.445 668.605 -14.115 ;
        RECT 666.915 -14.445 667.245 -14.115 ;
        RECT 665.555 -14.445 665.885 -14.115 ;
        RECT 664.195 -14.445 664.525 -14.115 ;
        RECT 662.835 -14.445 663.165 -14.115 ;
        RECT 661.475 -14.445 661.805 -14.115 ;
        RECT 660.115 -14.445 660.445 -14.115 ;
        RECT 658.755 -14.445 659.085 -14.115 ;
        RECT 657.395 -14.445 657.725 -14.115 ;
        RECT 656.035 -14.445 656.365 -14.115 ;
        RECT 654.675 -14.445 655.005 -14.115 ;
        RECT 653.315 -14.445 653.645 -14.115 ;
        RECT 651.955 -14.445 652.285 -14.115 ;
        RECT 650.595 -14.445 650.925 -14.115 ;
        RECT 649.235 -14.445 649.565 -14.115 ;
        RECT 647.875 -14.445 648.205 -14.115 ;
        RECT 646.515 -14.445 646.845 -14.115 ;
        RECT 645.155 -14.445 645.485 -14.115 ;
        RECT 643.795 -14.445 644.125 -14.115 ;
        RECT 642.435 -14.445 642.765 -14.115 ;
        RECT 641.075 -14.445 641.405 -14.115 ;
        RECT 639.715 -14.445 640.045 -14.115 ;
        RECT 638.355 -14.445 638.685 -14.115 ;
        RECT 636.995 -14.445 637.325 -14.115 ;
        RECT 635.635 -14.445 635.965 -14.115 ;
        RECT 634.275 -14.445 634.605 -14.115 ;
        RECT 632.915 -14.445 633.245 -14.115 ;
        RECT 631.555 -14.445 631.885 -14.115 ;
        RECT 630.195 -14.445 630.525 -14.115 ;
        RECT 628.835 -14.445 629.165 -14.115 ;
        RECT 627.475 -14.445 627.805 -14.115 ;
        RECT 626.115 -14.445 626.445 -14.115 ;
        RECT 624.755 -14.445 625.085 -14.115 ;
        RECT 623.395 -14.445 623.725 -14.115 ;
        RECT 622.035 -14.445 622.365 -14.115 ;
        RECT 620.675 -14.445 621.005 -14.115 ;
        RECT 619.315 -14.445 619.645 -14.115 ;
        RECT 617.955 -14.445 618.285 -14.115 ;
        RECT 616.595 -14.445 616.925 -14.115 ;
        RECT 615.235 -14.445 615.565 -14.115 ;
        RECT 613.875 -14.445 614.205 -14.115 ;
        RECT 612.515 -14.445 612.845 -14.115 ;
        RECT 611.155 -14.445 611.485 -14.115 ;
        RECT 609.795 -14.445 610.125 -14.115 ;
        RECT 608.435 -14.445 608.765 -14.115 ;
        RECT 607.075 -14.445 607.405 -14.115 ;
        RECT 605.715 -14.445 606.045 -14.115 ;
        RECT 604.355 -14.445 604.685 -14.115 ;
        RECT 602.995 -14.445 603.325 -14.115 ;
        RECT 601.635 -14.445 601.965 -14.115 ;
        RECT 600.275 -14.445 600.605 -14.115 ;
        RECT 598.915 -14.445 599.245 -14.115 ;
        RECT 597.555 -14.445 597.885 -14.115 ;
        RECT 596.195 -14.445 596.525 -14.115 ;
        RECT 594.835 -14.445 595.165 -14.115 ;
        RECT 593.475 -14.445 593.805 -14.115 ;
        RECT 592.115 -14.445 592.445 -14.115 ;
        RECT 590.755 -14.445 591.085 -14.115 ;
        RECT 589.395 -14.445 589.725 -14.115 ;
        RECT 588.035 -14.445 588.365 -14.115 ;
        RECT 586.675 -14.445 587.005 -14.115 ;
        RECT 585.315 -14.445 585.645 -14.115 ;
        RECT 583.955 -14.445 584.285 -14.115 ;
        RECT 582.595 -14.445 582.925 -14.115 ;
        RECT 581.235 -14.445 581.565 -14.115 ;
        RECT 579.875 -14.445 580.205 -14.115 ;
        RECT 578.515 -14.445 578.845 -14.115 ;
        RECT 577.155 -14.445 577.485 -14.115 ;
        RECT 575.795 -14.445 576.125 -14.115 ;
        RECT 574.435 -14.445 574.765 -14.115 ;
        RECT 573.075 -14.445 573.405 -14.115 ;
        RECT 571.715 -14.445 572.045 -14.115 ;
        RECT 570.355 -14.445 570.685 -14.115 ;
        RECT 568.995 -14.445 569.325 -14.115 ;
        RECT 567.635 -14.445 567.965 -14.115 ;
        RECT 566.275 -14.445 566.605 -14.115 ;
        RECT 564.915 -14.445 565.245 -14.115 ;
        RECT 563.555 -14.445 563.885 -14.115 ;
        RECT 562.195 -14.445 562.525 -14.115 ;
        RECT 560.835 -14.445 561.165 -14.115 ;
        RECT 559.475 -14.445 559.805 -14.115 ;
        RECT 558.115 -14.445 558.445 -14.115 ;
        RECT 556.755 -14.445 557.085 -14.115 ;
        RECT 555.395 -14.445 555.725 -14.115 ;
        RECT 554.035 -14.445 554.365 -14.115 ;
        RECT 552.675 -14.445 553.005 -14.115 ;
        RECT 551.315 -14.445 551.645 -14.115 ;
        RECT 549.955 -14.445 550.285 -14.115 ;
        RECT 548.595 -14.445 548.925 -14.115 ;
        RECT 547.235 -14.445 547.565 -14.115 ;
        RECT 545.875 -14.445 546.205 -14.115 ;
        RECT 544.515 -14.445 544.845 -14.115 ;
        RECT 543.155 -14.445 543.485 -14.115 ;
        RECT 541.795 -14.445 542.125 -14.115 ;
        RECT 540.435 -14.445 540.765 -14.115 ;
        RECT 539.075 -14.445 539.405 -14.115 ;
        RECT 537.715 -14.445 538.045 -14.115 ;
        RECT 536.355 -14.445 536.685 -14.115 ;
        RECT 534.995 -14.445 535.325 -14.115 ;
        RECT 533.635 -14.445 533.965 -14.115 ;
        RECT 532.275 -14.445 532.605 -14.115 ;
        RECT 530.915 -14.445 531.245 -14.115 ;
        RECT 529.555 -14.445 529.885 -14.115 ;
        RECT 528.195 -14.445 528.525 -14.115 ;
        RECT 526.835 -14.445 527.165 -14.115 ;
        RECT 525.475 -14.445 525.805 -14.115 ;
        RECT 524.115 -14.445 524.445 -14.115 ;
        RECT 522.755 -14.445 523.085 -14.115 ;
        RECT 521.395 -14.445 521.725 -14.115 ;
        RECT 520.035 -14.445 520.365 -14.115 ;
        RECT 518.675 -14.445 519.005 -14.115 ;
        RECT 517.315 -14.445 517.645 -14.115 ;
        RECT 515.955 -14.445 516.285 -14.115 ;
        RECT 514.595 -14.445 514.925 -14.115 ;
        RECT 513.235 -14.445 513.565 -14.115 ;
        RECT 511.875 -14.445 512.205 -14.115 ;
        RECT 510.515 -14.445 510.845 -14.115 ;
        RECT 509.155 -14.445 509.485 -14.115 ;
        RECT 507.795 -14.445 508.125 -14.115 ;
        RECT 506.435 -14.445 506.765 -14.115 ;
        RECT 505.075 -14.445 505.405 -14.115 ;
        RECT 503.715 -14.445 504.045 -14.115 ;
        RECT 502.355 -14.445 502.685 -14.115 ;
        RECT 500.995 -14.445 501.325 -14.115 ;
        RECT 499.635 -14.445 499.965 -14.115 ;
        RECT 498.275 -14.445 498.605 -14.115 ;
        RECT 496.915 -14.445 497.245 -14.115 ;
        RECT 495.555 -14.445 495.885 -14.115 ;
        RECT 494.195 -14.445 494.525 -14.115 ;
        RECT 492.835 -14.445 493.165 -14.115 ;
        RECT 491.475 -14.445 491.805 -14.115 ;
        RECT 490.115 -14.445 490.445 -14.115 ;
        RECT 488.755 -14.445 489.085 -14.115 ;
        RECT 487.395 -14.445 487.725 -14.115 ;
        RECT 486.035 -14.445 486.365 -14.115 ;
        RECT 484.675 -14.445 485.005 -14.115 ;
        RECT 483.315 -14.445 483.645 -14.115 ;
        RECT 481.955 -14.445 482.285 -14.115 ;
        RECT 480.595 -14.445 480.925 -14.115 ;
        RECT 479.235 -14.445 479.565 -14.115 ;
        RECT 477.875 -14.445 478.205 -14.115 ;
        RECT 476.515 -14.445 476.845 -14.115 ;
        RECT 475.155 -14.445 475.485 -14.115 ;
        RECT 473.795 -14.445 474.125 -14.115 ;
        RECT 472.435 -14.445 472.765 -14.115 ;
        RECT 471.075 -14.445 471.405 -14.115 ;
        RECT 469.715 -14.445 470.045 -14.115 ;
        RECT 468.355 -14.445 468.685 -14.115 ;
        RECT 466.995 -14.445 467.325 -14.115 ;
        RECT 465.635 -14.445 465.965 -14.115 ;
        RECT 464.275 -14.445 464.605 -14.115 ;
        RECT 462.915 -14.445 463.245 -14.115 ;
        RECT 461.555 -14.445 461.885 -14.115 ;
        RECT 460.195 -14.445 460.525 -14.115 ;
        RECT 458.835 -14.445 459.165 -14.115 ;
        RECT 457.475 -14.445 457.805 -14.115 ;
        RECT 456.115 -14.445 456.445 -14.115 ;
        RECT 454.755 -14.445 455.085 -14.115 ;
        RECT 453.395 -14.445 453.725 -14.115 ;
        RECT 452.035 -14.445 452.365 -14.115 ;
        RECT 450.675 -14.445 451.005 -14.115 ;
        RECT 449.315 -14.445 449.645 -14.115 ;
        RECT 447.955 -14.445 448.285 -14.115 ;
        RECT 446.595 -14.445 446.925 -14.115 ;
        RECT 445.235 -14.445 445.565 -14.115 ;
        RECT 443.875 -14.445 444.205 -14.115 ;
        RECT 442.515 -14.445 442.845 -14.115 ;
        RECT 441.155 -14.445 441.485 -14.115 ;
        RECT 439.795 -14.445 440.125 -14.115 ;
        RECT 438.435 -14.445 438.765 -14.115 ;
        RECT 437.075 -14.445 437.405 -14.115 ;
        RECT 435.715 -14.445 436.045 -14.115 ;
        RECT 434.355 -14.445 434.685 -14.115 ;
        RECT 432.995 -14.445 433.325 -14.115 ;
        RECT 431.635 -14.445 431.965 -14.115 ;
        RECT 430.275 -14.445 430.605 -14.115 ;
        RECT 428.915 -14.445 429.245 -14.115 ;
        RECT 427.555 -14.445 427.885 -14.115 ;
        RECT 426.195 -14.445 426.525 -14.115 ;
        RECT 424.835 -14.445 425.165 -14.115 ;
        RECT 423.475 -14.445 423.805 -14.115 ;
        RECT 422.115 -14.445 422.445 -14.115 ;
        RECT 420.755 -14.445 421.085 -14.115 ;
        RECT 419.395 -14.445 419.725 -14.115 ;
        RECT 418.035 -14.445 418.365 -14.115 ;
        RECT 416.675 -14.445 417.005 -14.115 ;
        RECT 415.315 -14.445 415.645 -14.115 ;
        RECT 413.955 -14.445 414.285 -14.115 ;
        RECT 412.595 -14.445 412.925 -14.115 ;
        RECT 411.235 -14.445 411.565 -14.115 ;
        RECT 409.875 -14.445 410.205 -14.115 ;
        RECT 408.515 -14.445 408.845 -14.115 ;
        RECT 407.155 -14.445 407.485 -14.115 ;
        RECT 405.795 -14.445 406.125 -14.115 ;
        RECT 404.435 -14.445 404.765 -14.115 ;
        RECT 403.075 -14.445 403.405 -14.115 ;
        RECT 401.715 -14.445 402.045 -14.115 ;
        RECT 400.355 -14.445 400.685 -14.115 ;
        RECT 398.995 -14.445 399.325 -14.115 ;
        RECT 397.635 -14.445 397.965 -14.115 ;
        RECT 396.275 -14.445 396.605 -14.115 ;
        RECT 394.915 -14.445 395.245 -14.115 ;
        RECT 393.555 -14.445 393.885 -14.115 ;
        RECT 392.195 -14.445 392.525 -14.115 ;
        RECT 390.835 -14.445 391.165 -14.115 ;
        RECT 389.475 -14.445 389.805 -14.115 ;
        RECT 388.115 -14.445 388.445 -14.115 ;
        RECT 386.755 -14.445 387.085 -14.115 ;
        RECT 385.395 -14.445 385.725 -14.115 ;
        RECT 384.035 -14.445 384.365 -14.115 ;
        RECT 382.675 -14.445 383.005 -14.115 ;
        RECT 381.315 -14.445 381.645 -14.115 ;
        RECT 379.955 -14.445 380.285 -14.115 ;
        RECT 378.595 -14.445 378.925 -14.115 ;
        RECT 377.235 -14.445 377.565 -14.115 ;
        RECT 375.875 -14.445 376.205 -14.115 ;
        RECT 374.515 -14.445 374.845 -14.115 ;
        RECT 373.155 -14.445 373.485 -14.115 ;
        RECT 371.795 -14.445 372.125 -14.115 ;
        RECT 370.435 -14.445 370.765 -14.115 ;
        RECT 369.075 -14.445 369.405 -14.115 ;
        RECT 367.715 -14.445 368.045 -14.115 ;
        RECT 366.355 -14.445 366.685 -14.115 ;
        RECT 364.995 -14.445 365.325 -14.115 ;
        RECT 363.635 -14.445 363.965 -14.115 ;
        RECT 362.275 -14.445 362.605 -14.115 ;
        RECT 360.915 -14.445 361.245 -14.115 ;
        RECT 359.555 -14.445 359.885 -14.115 ;
        RECT 358.195 -14.445 358.525 -14.115 ;
        RECT 356.835 -14.445 357.165 -14.115 ;
        RECT 355.475 -14.445 355.805 -14.115 ;
        RECT 354.115 -14.445 354.445 -14.115 ;
        RECT 352.755 -14.445 353.085 -14.115 ;
        RECT 351.395 -14.445 351.725 -14.115 ;
        RECT 350.035 -14.445 350.365 -14.115 ;
        RECT 348.675 -14.445 349.005 -14.115 ;
        RECT 347.315 -14.445 347.645 -14.115 ;
        RECT 345.955 -14.445 346.285 -14.115 ;
        RECT 344.595 -14.445 344.925 -14.115 ;
        RECT 343.235 -14.445 343.565 -14.115 ;
        RECT 341.875 -14.445 342.205 -14.115 ;
        RECT 340.515 -14.445 340.845 -14.115 ;
        RECT 339.155 -14.445 339.485 -14.115 ;
        RECT 337.795 -14.445 338.125 -14.115 ;
        RECT 336.435 -14.445 336.765 -14.115 ;
        RECT 335.075 -14.445 335.405 -14.115 ;
        RECT 333.715 -14.445 334.045 -14.115 ;
        RECT 332.355 -14.445 332.685 -14.115 ;
        RECT 330.995 -14.445 331.325 -14.115 ;
        RECT 329.635 -14.445 329.965 -14.115 ;
        RECT 328.275 -14.445 328.605 -14.115 ;
        RECT 326.915 -14.445 327.245 -14.115 ;
        RECT 325.555 -14.445 325.885 -14.115 ;
        RECT 324.195 -14.445 324.525 -14.115 ;
        RECT 322.835 -14.445 323.165 -14.115 ;
        RECT 321.475 -14.445 321.805 -14.115 ;
        RECT 320.115 -14.445 320.445 -14.115 ;
        RECT 318.755 -14.445 319.085 -14.115 ;
        RECT 317.395 -14.445 317.725 -14.115 ;
        RECT 316.035 -14.445 316.365 -14.115 ;
        RECT 314.675 -14.445 315.005 -14.115 ;
        RECT 313.315 -14.445 313.645 -14.115 ;
        RECT 311.955 -14.445 312.285 -14.115 ;
        RECT 310.595 -14.445 310.925 -14.115 ;
        RECT 309.235 -14.445 309.565 -14.115 ;
        RECT 307.875 -14.445 308.205 -14.115 ;
        RECT 306.515 -14.445 306.845 -14.115 ;
        RECT 305.155 -14.445 305.485 -14.115 ;
        RECT 303.795 -14.445 304.125 -14.115 ;
        RECT 302.435 -14.445 302.765 -14.115 ;
        RECT 301.075 -14.445 301.405 -14.115 ;
        RECT 299.715 -14.445 300.045 -14.115 ;
        RECT 298.355 -14.445 298.685 -14.115 ;
        RECT 296.995 -14.445 297.325 -14.115 ;
        RECT 295.635 -14.445 295.965 -14.115 ;
        RECT 294.275 -14.445 294.605 -14.115 ;
        RECT 292.915 -14.445 293.245 -14.115 ;
        RECT 291.555 -14.445 291.885 -14.115 ;
        RECT 290.195 -14.445 290.525 -14.115 ;
        RECT 288.835 -14.445 289.165 -14.115 ;
        RECT 287.475 -14.445 287.805 -14.115 ;
        RECT 286.115 -14.445 286.445 -14.115 ;
        RECT 284.755 -14.445 285.085 -14.115 ;
        RECT 283.395 -14.445 283.725 -14.115 ;
        RECT 282.035 -14.445 282.365 -14.115 ;
        RECT 280.675 -14.445 281.005 -14.115 ;
        RECT 279.315 -14.445 279.645 -14.115 ;
        RECT 277.955 -14.445 278.285 -14.115 ;
        RECT 276.595 -14.445 276.925 -14.115 ;
        RECT 275.235 -14.445 275.565 -14.115 ;
        RECT 273.875 -14.445 274.205 -14.115 ;
        RECT 272.515 -14.445 272.845 -14.115 ;
        RECT 271.155 -14.445 271.485 -14.115 ;
        RECT 269.795 -14.445 270.125 -14.115 ;
        RECT 268.435 -14.445 268.765 -14.115 ;
        RECT 267.075 -14.445 267.405 -14.115 ;
        RECT 265.715 -14.445 266.045 -14.115 ;
        RECT 264.355 -14.445 264.685 -14.115 ;
        RECT 262.995 -14.445 263.325 -14.115 ;
        RECT 261.635 -14.445 261.965 -14.115 ;
        RECT 260.275 -14.445 260.605 -14.115 ;
        RECT 258.915 -14.445 259.245 -14.115 ;
        RECT 257.555 -14.445 257.885 -14.115 ;
        RECT 256.195 -14.445 256.525 -14.115 ;
        RECT 254.835 -14.445 255.165 -14.115 ;
        RECT 253.475 -14.445 253.805 -14.115 ;
        RECT 252.115 -14.445 252.445 -14.115 ;
        RECT 250.755 -14.445 251.085 -14.115 ;
        RECT 249.395 -14.445 249.725 -14.115 ;
        RECT 248.035 -14.445 248.365 -14.115 ;
        RECT 246.675 -14.445 247.005 -14.115 ;
        RECT 245.315 -14.445 245.645 -14.115 ;
        RECT 243.955 -14.445 244.285 -14.115 ;
        RECT 242.595 -14.445 242.925 -14.115 ;
        RECT 241.235 -14.445 241.565 -14.115 ;
        RECT 239.875 -14.445 240.205 -14.115 ;
        RECT 238.515 -14.445 238.845 -14.115 ;
        RECT 237.155 -14.445 237.485 -14.115 ;
        RECT 235.795 -14.445 236.125 -14.115 ;
        RECT 234.435 -14.445 234.765 -14.115 ;
        RECT 233.075 -14.445 233.405 -14.115 ;
        RECT 231.715 -14.445 232.045 -14.115 ;
        RECT 230.355 -14.445 230.685 -14.115 ;
        RECT 228.995 -14.445 229.325 -14.115 ;
        RECT 227.635 -14.445 227.965 -14.115 ;
        RECT 226.275 -14.445 226.605 -14.115 ;
        RECT 224.915 -14.445 225.245 -14.115 ;
        RECT 223.555 -14.445 223.885 -14.115 ;
        RECT 222.195 -14.445 222.525 -14.115 ;
        RECT 220.835 -14.445 221.165 -14.115 ;
        RECT 219.475 -14.445 219.805 -14.115 ;
        RECT 218.115 -14.445 218.445 -14.115 ;
        RECT 216.755 -14.445 217.085 -14.115 ;
        RECT 215.395 -14.445 215.725 -14.115 ;
        RECT 214.035 -14.445 214.365 -14.115 ;
        RECT 212.675 -14.445 213.005 -14.115 ;
        RECT 211.315 -14.445 211.645 -14.115 ;
        RECT 209.955 -14.445 210.285 -14.115 ;
        RECT 208.595 -14.445 208.925 -14.115 ;
        RECT 207.235 -14.445 207.565 -14.115 ;
        RECT 205.875 -14.445 206.205 -14.115 ;
        RECT 204.515 -14.445 204.845 -14.115 ;
        RECT 203.155 -14.445 203.485 -14.115 ;
        RECT 201.795 -14.445 202.125 -14.115 ;
        RECT 200.435 -14.445 200.765 -14.115 ;
        RECT 199.075 -14.445 199.405 -14.115 ;
        RECT 197.715 -14.445 198.045 -14.115 ;
        RECT 196.355 -14.445 196.685 -14.115 ;
        RECT 194.995 -14.445 195.325 -14.115 ;
        RECT 193.635 -14.445 193.965 -14.115 ;
        RECT 192.275 -14.445 192.605 -14.115 ;
        RECT 190.915 -14.445 191.245 -14.115 ;
        RECT 189.555 -14.445 189.885 -14.115 ;
        RECT 188.195 -14.445 188.525 -14.115 ;
        RECT 186.835 -14.445 187.165 -14.115 ;
        RECT 185.475 -14.445 185.805 -14.115 ;
        RECT 184.115 -14.445 184.445 -14.115 ;
        RECT 182.755 -14.445 183.085 -14.115 ;
        RECT 181.395 -14.445 181.725 -14.115 ;
        RECT 180.035 -14.445 180.365 -14.115 ;
        RECT 178.675 -14.445 179.005 -14.115 ;
        RECT 177.315 -14.445 177.645 -14.115 ;
        RECT 175.955 -14.445 176.285 -14.115 ;
        RECT 174.595 -14.445 174.925 -14.115 ;
        RECT 173.235 -14.445 173.565 -14.115 ;
        RECT 171.875 -14.445 172.205 -14.115 ;
        RECT 170.515 -14.445 170.845 -14.115 ;
        RECT 169.155 -14.445 169.485 -14.115 ;
        RECT 167.795 -14.445 168.125 -14.115 ;
        RECT 166.435 -14.445 166.765 -14.115 ;
        RECT 165.075 -14.445 165.405 -14.115 ;
        RECT 163.715 -14.445 164.045 -14.115 ;
        RECT 162.355 -14.445 162.685 -14.115 ;
        RECT 160.995 -14.445 161.325 -14.115 ;
        RECT 159.635 -14.445 159.965 -14.115 ;
        RECT 158.275 -14.445 158.605 -14.115 ;
        RECT 156.915 -14.445 157.245 -14.115 ;
        RECT 155.555 -14.445 155.885 -14.115 ;
        RECT 154.195 -14.445 154.525 -14.115 ;
        RECT 152.835 -14.445 153.165 -14.115 ;
        RECT 151.475 -14.445 151.805 -14.115 ;
        RECT 150.115 -14.445 150.445 -14.115 ;
        RECT 148.755 -14.445 149.085 -14.115 ;
        RECT 147.395 -14.445 147.725 -14.115 ;
        RECT 146.035 -14.445 146.365 -14.115 ;
        RECT 144.675 -14.445 145.005 -14.115 ;
        RECT 143.315 -14.445 143.645 -14.115 ;
        RECT 141.955 -14.445 142.285 -14.115 ;
        RECT 140.595 -14.445 140.925 -14.115 ;
        RECT 139.235 -14.445 139.565 -14.115 ;
        RECT 137.875 -14.445 138.205 -14.115 ;
        RECT 136.515 -14.445 136.845 -14.115 ;
        RECT 135.155 -14.445 135.485 -14.115 ;
        RECT 133.795 -14.445 134.125 -14.115 ;
        RECT 132.435 -14.445 132.765 -14.115 ;
        RECT 131.075 -14.445 131.405 -14.115 ;
        RECT 129.715 -14.445 130.045 -14.115 ;
        RECT 128.355 -14.445 128.685 -14.115 ;
        RECT 126.995 -14.445 127.325 -14.115 ;
        RECT 678.125 -14.44 954.88 -14.12 ;
        RECT 953.875 -14.445 954.205 -14.115 ;
        RECT 952.515 -14.445 952.845 -14.115 ;
        RECT 951.155 -14.445 951.485 -14.115 ;
        RECT 949.795 -14.445 950.125 -14.115 ;
        RECT 948.435 -14.445 948.765 -14.115 ;
        RECT 947.075 -14.445 947.405 -14.115 ;
        RECT 945.715 -14.445 946.045 -14.115 ;
        RECT 944.355 -14.445 944.685 -14.115 ;
        RECT 942.995 -14.445 943.325 -14.115 ;
        RECT 941.635 -14.445 941.965 -14.115 ;
        RECT 940.275 -14.445 940.605 -14.115 ;
        RECT 938.915 -14.445 939.245 -14.115 ;
        RECT 937.555 -14.445 937.885 -14.115 ;
        RECT 936.195 -14.445 936.525 -14.115 ;
        RECT 934.835 -14.445 935.165 -14.115 ;
        RECT 933.475 -14.445 933.805 -14.115 ;
        RECT 932.115 -14.445 932.445 -14.115 ;
        RECT 930.755 -14.445 931.085 -14.115 ;
        RECT 929.395 -14.445 929.725 -14.115 ;
        RECT 928.035 -14.445 928.365 -14.115 ;
        RECT 926.675 -14.445 927.005 -14.115 ;
        RECT 925.315 -14.445 925.645 -14.115 ;
        RECT 923.955 -14.445 924.285 -14.115 ;
        RECT 922.595 -14.445 922.925 -14.115 ;
        RECT 921.235 -14.445 921.565 -14.115 ;
        RECT 919.875 -14.445 920.205 -14.115 ;
        RECT 918.515 -14.445 918.845 -14.115 ;
        RECT 917.155 -14.445 917.485 -14.115 ;
        RECT 915.795 -14.445 916.125 -14.115 ;
        RECT 914.435 -14.445 914.765 -14.115 ;
        RECT 913.075 -14.445 913.405 -14.115 ;
        RECT 911.715 -14.445 912.045 -14.115 ;
        RECT 910.355 -14.445 910.685 -14.115 ;
        RECT 908.995 -14.445 909.325 -14.115 ;
        RECT 907.635 -14.445 907.965 -14.115 ;
        RECT 906.275 -14.445 906.605 -14.115 ;
        RECT 904.915 -14.445 905.245 -14.115 ;
        RECT 903.555 -14.445 903.885 -14.115 ;
        RECT 902.195 -14.445 902.525 -14.115 ;
        RECT 900.835 -14.445 901.165 -14.115 ;
        RECT 899.475 -14.445 899.805 -14.115 ;
        RECT 898.115 -14.445 898.445 -14.115 ;
        RECT 896.755 -14.445 897.085 -14.115 ;
        RECT 895.395 -14.445 895.725 -14.115 ;
        RECT 894.035 -14.445 894.365 -14.115 ;
        RECT 892.675 -14.445 893.005 -14.115 ;
        RECT 891.315 -14.445 891.645 -14.115 ;
        RECT 889.955 -14.445 890.285 -14.115 ;
        RECT 888.595 -14.445 888.925 -14.115 ;
        RECT 887.235 -14.445 887.565 -14.115 ;
        RECT 885.875 -14.445 886.205 -14.115 ;
        RECT 884.515 -14.445 884.845 -14.115 ;
        RECT 883.155 -14.445 883.485 -14.115 ;
        RECT 881.795 -14.445 882.125 -14.115 ;
        RECT 880.435 -14.445 880.765 -14.115 ;
        RECT 879.075 -14.445 879.405 -14.115 ;
        RECT 877.715 -14.445 878.045 -14.115 ;
        RECT 876.355 -14.445 876.685 -14.115 ;
        RECT 874.995 -14.445 875.325 -14.115 ;
        RECT 873.635 -14.445 873.965 -14.115 ;
        RECT 872.275 -14.445 872.605 -14.115 ;
        RECT 870.915 -14.445 871.245 -14.115 ;
        RECT 869.555 -14.445 869.885 -14.115 ;
        RECT 868.195 -14.445 868.525 -14.115 ;
        RECT 866.835 -14.445 867.165 -14.115 ;
        RECT 865.475 -14.445 865.805 -14.115 ;
        RECT 864.115 -14.445 864.445 -14.115 ;
        RECT 862.755 -14.445 863.085 -14.115 ;
        RECT 861.395 -14.445 861.725 -14.115 ;
        RECT 860.035 -14.445 860.365 -14.115 ;
        RECT 858.675 -14.445 859.005 -14.115 ;
        RECT 857.315 -14.445 857.645 -14.115 ;
        RECT 855.955 -14.445 856.285 -14.115 ;
        RECT 854.595 -14.445 854.925 -14.115 ;
        RECT 853.235 -14.445 853.565 -14.115 ;
        RECT 851.875 -14.445 852.205 -14.115 ;
        RECT 850.515 -14.445 850.845 -14.115 ;
        RECT 849.155 -14.445 849.485 -14.115 ;
        RECT 847.795 -14.445 848.125 -14.115 ;
        RECT 846.435 -14.445 846.765 -14.115 ;
        RECT 845.075 -14.445 845.405 -14.115 ;
        RECT 843.715 -14.445 844.045 -14.115 ;
        RECT 842.355 -14.445 842.685 -14.115 ;
        RECT 840.995 -14.445 841.325 -14.115 ;
        RECT 839.635 -14.445 839.965 -14.115 ;
        RECT 838.275 -14.445 838.605 -14.115 ;
        RECT 836.915 -14.445 837.245 -14.115 ;
        RECT 835.555 -14.445 835.885 -14.115 ;
        RECT 834.195 -14.445 834.525 -14.115 ;
        RECT 832.835 -14.445 833.165 -14.115 ;
        RECT 831.475 -14.445 831.805 -14.115 ;
        RECT 830.115 -14.445 830.445 -14.115 ;
        RECT 828.755 -14.445 829.085 -14.115 ;
        RECT 827.395 -14.445 827.725 -14.115 ;
        RECT 826.035 -14.445 826.365 -14.115 ;
        RECT 824.675 -14.445 825.005 -14.115 ;
        RECT 823.315 -14.445 823.645 -14.115 ;
        RECT 821.955 -14.445 822.285 -14.115 ;
        RECT 820.595 -14.445 820.925 -14.115 ;
        RECT 819.235 -14.445 819.565 -14.115 ;
        RECT 817.875 -14.445 818.205 -14.115 ;
        RECT 816.515 -14.445 816.845 -14.115 ;
        RECT 815.155 -14.445 815.485 -14.115 ;
        RECT 813.795 -14.445 814.125 -14.115 ;
        RECT 812.435 -14.445 812.765 -14.115 ;
        RECT 811.075 -14.445 811.405 -14.115 ;
        RECT 809.715 -14.445 810.045 -14.115 ;
        RECT 808.355 -14.445 808.685 -14.115 ;
        RECT 806.995 -14.445 807.325 -14.115 ;
        RECT 805.635 -14.445 805.965 -14.115 ;
        RECT 804.275 -14.445 804.605 -14.115 ;
        RECT 802.915 -14.445 803.245 -14.115 ;
        RECT 801.555 -14.445 801.885 -14.115 ;
        RECT 800.195 -14.445 800.525 -14.115 ;
        RECT 798.835 -14.445 799.165 -14.115 ;
        RECT 797.475 -14.445 797.805 -14.115 ;
        RECT 796.115 -14.445 796.445 -14.115 ;
        RECT 794.755 -14.445 795.085 -14.115 ;
        RECT 793.395 -14.445 793.725 -14.115 ;
        RECT 792.035 -14.445 792.365 -14.115 ;
        RECT 790.675 -14.445 791.005 -14.115 ;
        RECT 789.315 -14.445 789.645 -14.115 ;
        RECT 787.955 -14.445 788.285 -14.115 ;
        RECT 786.595 -14.445 786.925 -14.115 ;
        RECT 785.235 -14.445 785.565 -14.115 ;
        RECT 783.875 -14.445 784.205 -14.115 ;
        RECT 782.515 -14.445 782.845 -14.115 ;
        RECT 781.155 -14.445 781.485 -14.115 ;
        RECT 779.795 -14.445 780.125 -14.115 ;
        RECT 778.435 -14.445 778.765 -14.115 ;
        RECT 777.075 -14.445 777.405 -14.115 ;
        RECT 775.715 -14.445 776.045 -14.115 ;
        RECT 774.355 -14.445 774.685 -14.115 ;
        RECT 772.995 -14.445 773.325 -14.115 ;
        RECT 771.635 -14.445 771.965 -14.115 ;
        RECT 770.275 -14.445 770.605 -14.115 ;
        RECT 768.915 -14.445 769.245 -14.115 ;
        RECT 767.555 -14.445 767.885 -14.115 ;
        RECT 766.195 -14.445 766.525 -14.115 ;
        RECT 764.835 -14.445 765.165 -14.115 ;
        RECT 763.475 -14.445 763.805 -14.115 ;
        RECT 762.115 -14.445 762.445 -14.115 ;
        RECT 760.755 -14.445 761.085 -14.115 ;
        RECT 759.395 -14.445 759.725 -14.115 ;
        RECT 758.035 -14.445 758.365 -14.115 ;
        RECT 756.675 -14.445 757.005 -14.115 ;
        RECT 755.315 -14.445 755.645 -14.115 ;
        RECT 753.955 -14.445 754.285 -14.115 ;
        RECT 752.595 -14.445 752.925 -14.115 ;
        RECT 751.235 -14.445 751.565 -14.115 ;
        RECT 749.875 -14.445 750.205 -14.115 ;
        RECT 748.515 -14.445 748.845 -14.115 ;
        RECT 747.155 -14.445 747.485 -14.115 ;
        RECT 745.795 -14.445 746.125 -14.115 ;
        RECT 744.435 -14.445 744.765 -14.115 ;
        RECT 743.075 -14.445 743.405 -14.115 ;
        RECT 741.715 -14.445 742.045 -14.115 ;
        RECT 740.355 -14.445 740.685 -14.115 ;
        RECT 738.995 -14.445 739.325 -14.115 ;
        RECT 737.635 -14.445 737.965 -14.115 ;
        RECT 736.275 -14.445 736.605 -14.115 ;
        RECT 734.915 -14.445 735.245 -14.115 ;
        RECT 733.555 -14.445 733.885 -14.115 ;
        RECT 732.195 -14.445 732.525 -14.115 ;
        RECT 730.835 -14.445 731.165 -14.115 ;
        RECT 729.475 -14.445 729.805 -14.115 ;
        RECT 728.115 -14.445 728.445 -14.115 ;
        RECT 726.755 -14.445 727.085 -14.115 ;
        RECT 725.395 -14.445 725.725 -14.115 ;
        RECT 724.035 -14.445 724.365 -14.115 ;
        RECT 722.675 -14.445 723.005 -14.115 ;
        RECT 721.315 -14.445 721.645 -14.115 ;
        RECT 719.955 -14.445 720.285 -14.115 ;
        RECT 718.595 -14.445 718.925 -14.115 ;
        RECT 717.235 -14.445 717.565 -14.115 ;
        RECT 715.875 -14.445 716.205 -14.115 ;
        RECT 714.515 -14.445 714.845 -14.115 ;
        RECT 713.155 -14.445 713.485 -14.115 ;
        RECT 711.795 -14.445 712.125 -14.115 ;
        RECT 710.435 -14.445 710.765 -14.115 ;
        RECT 709.075 -14.445 709.405 -14.115 ;
        RECT 707.715 -14.445 708.045 -14.115 ;
        RECT 706.355 -14.445 706.685 -14.115 ;
        RECT 704.995 -14.445 705.325 -14.115 ;
        RECT 703.635 -14.445 703.965 -14.115 ;
        RECT 702.275 -14.445 702.605 -14.115 ;
        RECT 700.915 -14.445 701.245 -14.115 ;
        RECT 699.555 -14.445 699.885 -14.115 ;
        RECT 698.195 -14.445 698.525 -14.115 ;
        RECT 696.835 -14.445 697.165 -14.115 ;
        RECT 695.475 -14.445 695.805 -14.115 ;
        RECT 694.115 -14.445 694.445 -14.115 ;
        RECT 692.755 -14.445 693.085 -14.115 ;
        RECT 691.395 -14.445 691.725 -14.115 ;
        RECT 690.035 -14.445 690.365 -14.115 ;
        RECT 688.675 -14.445 689.005 -14.115 ;
        RECT 687.315 -14.445 687.645 -14.115 ;
        RECT 685.955 -14.445 686.285 -14.115 ;
        RECT 684.595 -14.445 684.925 -14.115 ;
        RECT 683.235 -14.445 683.565 -14.115 ;
        RECT 681.875 -14.445 682.205 -14.115 ;
        RECT 680.515 -14.445 680.845 -14.115 ;
        RECT 679.155 -14.445 679.485 -14.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 -10.365 678.125 -10.035 ;
        RECT -1.52 -10.36 678.125 -10.04 ;
        RECT 676.435 -10.365 676.765 -10.035 ;
        RECT 675.075 -10.365 675.405 -10.035 ;
        RECT 673.715 -10.365 674.045 -10.035 ;
        RECT 672.355 -10.365 672.685 -10.035 ;
        RECT 670.995 -10.365 671.325 -10.035 ;
        RECT 669.635 -10.365 669.965 -10.035 ;
        RECT 668.275 -10.365 668.605 -10.035 ;
        RECT 666.915 -10.365 667.245 -10.035 ;
        RECT 665.555 -10.365 665.885 -10.035 ;
        RECT 664.195 -10.365 664.525 -10.035 ;
        RECT 662.835 -10.365 663.165 -10.035 ;
        RECT 661.475 -10.365 661.805 -10.035 ;
        RECT 660.115 -10.365 660.445 -10.035 ;
        RECT 658.755 -10.365 659.085 -10.035 ;
        RECT 657.395 -10.365 657.725 -10.035 ;
        RECT 656.035 -10.365 656.365 -10.035 ;
        RECT 654.675 -10.365 655.005 -10.035 ;
        RECT 653.315 -10.365 653.645 -10.035 ;
        RECT 651.955 -10.365 652.285 -10.035 ;
        RECT 650.595 -10.365 650.925 -10.035 ;
        RECT 649.235 -10.365 649.565 -10.035 ;
        RECT 647.875 -10.365 648.205 -10.035 ;
        RECT 646.515 -10.365 646.845 -10.035 ;
        RECT 645.155 -10.365 645.485 -10.035 ;
        RECT 643.795 -10.365 644.125 -10.035 ;
        RECT 642.435 -10.365 642.765 -10.035 ;
        RECT 641.075 -10.365 641.405 -10.035 ;
        RECT 639.715 -10.365 640.045 -10.035 ;
        RECT 638.355 -10.365 638.685 -10.035 ;
        RECT 636.995 -10.365 637.325 -10.035 ;
        RECT 635.635 -10.365 635.965 -10.035 ;
        RECT 634.275 -10.365 634.605 -10.035 ;
        RECT 632.915 -10.365 633.245 -10.035 ;
        RECT 631.555 -10.365 631.885 -10.035 ;
        RECT 630.195 -10.365 630.525 -10.035 ;
        RECT 628.835 -10.365 629.165 -10.035 ;
        RECT 627.475 -10.365 627.805 -10.035 ;
        RECT 626.115 -10.365 626.445 -10.035 ;
        RECT 624.755 -10.365 625.085 -10.035 ;
        RECT 623.395 -10.365 623.725 -10.035 ;
        RECT 622.035 -10.365 622.365 -10.035 ;
        RECT 620.675 -10.365 621.005 -10.035 ;
        RECT 619.315 -10.365 619.645 -10.035 ;
        RECT 617.955 -10.365 618.285 -10.035 ;
        RECT 616.595 -10.365 616.925 -10.035 ;
        RECT 615.235 -10.365 615.565 -10.035 ;
        RECT 613.875 -10.365 614.205 -10.035 ;
        RECT 612.515 -10.365 612.845 -10.035 ;
        RECT 611.155 -10.365 611.485 -10.035 ;
        RECT 609.795 -10.365 610.125 -10.035 ;
        RECT 608.435 -10.365 608.765 -10.035 ;
        RECT 607.075 -10.365 607.405 -10.035 ;
        RECT 605.715 -10.365 606.045 -10.035 ;
        RECT 604.355 -10.365 604.685 -10.035 ;
        RECT 602.995 -10.365 603.325 -10.035 ;
        RECT 601.635 -10.365 601.965 -10.035 ;
        RECT 600.275 -10.365 600.605 -10.035 ;
        RECT 598.915 -10.365 599.245 -10.035 ;
        RECT 597.555 -10.365 597.885 -10.035 ;
        RECT 596.195 -10.365 596.525 -10.035 ;
        RECT 594.835 -10.365 595.165 -10.035 ;
        RECT 593.475 -10.365 593.805 -10.035 ;
        RECT 592.115 -10.365 592.445 -10.035 ;
        RECT 590.755 -10.365 591.085 -10.035 ;
        RECT 589.395 -10.365 589.725 -10.035 ;
        RECT 588.035 -10.365 588.365 -10.035 ;
        RECT 586.675 -10.365 587.005 -10.035 ;
        RECT 585.315 -10.365 585.645 -10.035 ;
        RECT 583.955 -10.365 584.285 -10.035 ;
        RECT 582.595 -10.365 582.925 -10.035 ;
        RECT 581.235 -10.365 581.565 -10.035 ;
        RECT 579.875 -10.365 580.205 -10.035 ;
        RECT 578.515 -10.365 578.845 -10.035 ;
        RECT 577.155 -10.365 577.485 -10.035 ;
        RECT 575.795 -10.365 576.125 -10.035 ;
        RECT 574.435 -10.365 574.765 -10.035 ;
        RECT 573.075 -10.365 573.405 -10.035 ;
        RECT 571.715 -10.365 572.045 -10.035 ;
        RECT 570.355 -10.365 570.685 -10.035 ;
        RECT 568.995 -10.365 569.325 -10.035 ;
        RECT 567.635 -10.365 567.965 -10.035 ;
        RECT 566.275 -10.365 566.605 -10.035 ;
        RECT 564.915 -10.365 565.245 -10.035 ;
        RECT 563.555 -10.365 563.885 -10.035 ;
        RECT 562.195 -10.365 562.525 -10.035 ;
        RECT 560.835 -10.365 561.165 -10.035 ;
        RECT 559.475 -10.365 559.805 -10.035 ;
        RECT 558.115 -10.365 558.445 -10.035 ;
        RECT 556.755 -10.365 557.085 -10.035 ;
        RECT 555.395 -10.365 555.725 -10.035 ;
        RECT 554.035 -10.365 554.365 -10.035 ;
        RECT 552.675 -10.365 553.005 -10.035 ;
        RECT 551.315 -10.365 551.645 -10.035 ;
        RECT 549.955 -10.365 550.285 -10.035 ;
        RECT 548.595 -10.365 548.925 -10.035 ;
        RECT 547.235 -10.365 547.565 -10.035 ;
        RECT 545.875 -10.365 546.205 -10.035 ;
        RECT 544.515 -10.365 544.845 -10.035 ;
        RECT 543.155 -10.365 543.485 -10.035 ;
        RECT 541.795 -10.365 542.125 -10.035 ;
        RECT 540.435 -10.365 540.765 -10.035 ;
        RECT 539.075 -10.365 539.405 -10.035 ;
        RECT 537.715 -10.365 538.045 -10.035 ;
        RECT 536.355 -10.365 536.685 -10.035 ;
        RECT 534.995 -10.365 535.325 -10.035 ;
        RECT 533.635 -10.365 533.965 -10.035 ;
        RECT 532.275 -10.365 532.605 -10.035 ;
        RECT 530.915 -10.365 531.245 -10.035 ;
        RECT 529.555 -10.365 529.885 -10.035 ;
        RECT 528.195 -10.365 528.525 -10.035 ;
        RECT 526.835 -10.365 527.165 -10.035 ;
        RECT 525.475 -10.365 525.805 -10.035 ;
        RECT 524.115 -10.365 524.445 -10.035 ;
        RECT 522.755 -10.365 523.085 -10.035 ;
        RECT 521.395 -10.365 521.725 -10.035 ;
        RECT 520.035 -10.365 520.365 -10.035 ;
        RECT 518.675 -10.365 519.005 -10.035 ;
        RECT 517.315 -10.365 517.645 -10.035 ;
        RECT 515.955 -10.365 516.285 -10.035 ;
        RECT 514.595 -10.365 514.925 -10.035 ;
        RECT 513.235 -10.365 513.565 -10.035 ;
        RECT 511.875 -10.365 512.205 -10.035 ;
        RECT 510.515 -10.365 510.845 -10.035 ;
        RECT 509.155 -10.365 509.485 -10.035 ;
        RECT 507.795 -10.365 508.125 -10.035 ;
        RECT 506.435 -10.365 506.765 -10.035 ;
        RECT 505.075 -10.365 505.405 -10.035 ;
        RECT 503.715 -10.365 504.045 -10.035 ;
        RECT 502.355 -10.365 502.685 -10.035 ;
        RECT 500.995 -10.365 501.325 -10.035 ;
        RECT 499.635 -10.365 499.965 -10.035 ;
        RECT 498.275 -10.365 498.605 -10.035 ;
        RECT 496.915 -10.365 497.245 -10.035 ;
        RECT 495.555 -10.365 495.885 -10.035 ;
        RECT 494.195 -10.365 494.525 -10.035 ;
        RECT 492.835 -10.365 493.165 -10.035 ;
        RECT 491.475 -10.365 491.805 -10.035 ;
        RECT 490.115 -10.365 490.445 -10.035 ;
        RECT 488.755 -10.365 489.085 -10.035 ;
        RECT 487.395 -10.365 487.725 -10.035 ;
        RECT 486.035 -10.365 486.365 -10.035 ;
        RECT 484.675 -10.365 485.005 -10.035 ;
        RECT 483.315 -10.365 483.645 -10.035 ;
        RECT 481.955 -10.365 482.285 -10.035 ;
        RECT 480.595 -10.365 480.925 -10.035 ;
        RECT 479.235 -10.365 479.565 -10.035 ;
        RECT 477.875 -10.365 478.205 -10.035 ;
        RECT 476.515 -10.365 476.845 -10.035 ;
        RECT 475.155 -10.365 475.485 -10.035 ;
        RECT 473.795 -10.365 474.125 -10.035 ;
        RECT 472.435 -10.365 472.765 -10.035 ;
        RECT 471.075 -10.365 471.405 -10.035 ;
        RECT 469.715 -10.365 470.045 -10.035 ;
        RECT 468.355 -10.365 468.685 -10.035 ;
        RECT 466.995 -10.365 467.325 -10.035 ;
        RECT 465.635 -10.365 465.965 -10.035 ;
        RECT 464.275 -10.365 464.605 -10.035 ;
        RECT 462.915 -10.365 463.245 -10.035 ;
        RECT 461.555 -10.365 461.885 -10.035 ;
        RECT 460.195 -10.365 460.525 -10.035 ;
        RECT 458.835 -10.365 459.165 -10.035 ;
        RECT 457.475 -10.365 457.805 -10.035 ;
        RECT 456.115 -10.365 456.445 -10.035 ;
        RECT 454.755 -10.365 455.085 -10.035 ;
        RECT 453.395 -10.365 453.725 -10.035 ;
        RECT 452.035 -10.365 452.365 -10.035 ;
        RECT 450.675 -10.365 451.005 -10.035 ;
        RECT 449.315 -10.365 449.645 -10.035 ;
        RECT 447.955 -10.365 448.285 -10.035 ;
        RECT 446.595 -10.365 446.925 -10.035 ;
        RECT 445.235 -10.365 445.565 -10.035 ;
        RECT 443.875 -10.365 444.205 -10.035 ;
        RECT 442.515 -10.365 442.845 -10.035 ;
        RECT 441.155 -10.365 441.485 -10.035 ;
        RECT 439.795 -10.365 440.125 -10.035 ;
        RECT 438.435 -10.365 438.765 -10.035 ;
        RECT 437.075 -10.365 437.405 -10.035 ;
        RECT 435.715 -10.365 436.045 -10.035 ;
        RECT 434.355 -10.365 434.685 -10.035 ;
        RECT 432.995 -10.365 433.325 -10.035 ;
        RECT 431.635 -10.365 431.965 -10.035 ;
        RECT 430.275 -10.365 430.605 -10.035 ;
        RECT 428.915 -10.365 429.245 -10.035 ;
        RECT 427.555 -10.365 427.885 -10.035 ;
        RECT 426.195 -10.365 426.525 -10.035 ;
        RECT 424.835 -10.365 425.165 -10.035 ;
        RECT 423.475 -10.365 423.805 -10.035 ;
        RECT 422.115 -10.365 422.445 -10.035 ;
        RECT 420.755 -10.365 421.085 -10.035 ;
        RECT 419.395 -10.365 419.725 -10.035 ;
        RECT 418.035 -10.365 418.365 -10.035 ;
        RECT 416.675 -10.365 417.005 -10.035 ;
        RECT 415.315 -10.365 415.645 -10.035 ;
        RECT 413.955 -10.365 414.285 -10.035 ;
        RECT 412.595 -10.365 412.925 -10.035 ;
        RECT 411.235 -10.365 411.565 -10.035 ;
        RECT 409.875 -10.365 410.205 -10.035 ;
        RECT 408.515 -10.365 408.845 -10.035 ;
        RECT 407.155 -10.365 407.485 -10.035 ;
        RECT 405.795 -10.365 406.125 -10.035 ;
        RECT 404.435 -10.365 404.765 -10.035 ;
        RECT 403.075 -10.365 403.405 -10.035 ;
        RECT 401.715 -10.365 402.045 -10.035 ;
        RECT 400.355 -10.365 400.685 -10.035 ;
        RECT 398.995 -10.365 399.325 -10.035 ;
        RECT 397.635 -10.365 397.965 -10.035 ;
        RECT 396.275 -10.365 396.605 -10.035 ;
        RECT 394.915 -10.365 395.245 -10.035 ;
        RECT 393.555 -10.365 393.885 -10.035 ;
        RECT 392.195 -10.365 392.525 -10.035 ;
        RECT 390.835 -10.365 391.165 -10.035 ;
        RECT 389.475 -10.365 389.805 -10.035 ;
        RECT 388.115 -10.365 388.445 -10.035 ;
        RECT 386.755 -10.365 387.085 -10.035 ;
        RECT 385.395 -10.365 385.725 -10.035 ;
        RECT 384.035 -10.365 384.365 -10.035 ;
        RECT 382.675 -10.365 383.005 -10.035 ;
        RECT 381.315 -10.365 381.645 -10.035 ;
        RECT 379.955 -10.365 380.285 -10.035 ;
        RECT 378.595 -10.365 378.925 -10.035 ;
        RECT 377.235 -10.365 377.565 -10.035 ;
        RECT 375.875 -10.365 376.205 -10.035 ;
        RECT 374.515 -10.365 374.845 -10.035 ;
        RECT 373.155 -10.365 373.485 -10.035 ;
        RECT 371.795 -10.365 372.125 -10.035 ;
        RECT 370.435 -10.365 370.765 -10.035 ;
        RECT 369.075 -10.365 369.405 -10.035 ;
        RECT 367.715 -10.365 368.045 -10.035 ;
        RECT 366.355 -10.365 366.685 -10.035 ;
        RECT 364.995 -10.365 365.325 -10.035 ;
        RECT 363.635 -10.365 363.965 -10.035 ;
        RECT 362.275 -10.365 362.605 -10.035 ;
        RECT 360.915 -10.365 361.245 -10.035 ;
        RECT 359.555 -10.365 359.885 -10.035 ;
        RECT 358.195 -10.365 358.525 -10.035 ;
        RECT 356.835 -10.365 357.165 -10.035 ;
        RECT 355.475 -10.365 355.805 -10.035 ;
        RECT 354.115 -10.365 354.445 -10.035 ;
        RECT 352.755 -10.365 353.085 -10.035 ;
        RECT 351.395 -10.365 351.725 -10.035 ;
        RECT 350.035 -10.365 350.365 -10.035 ;
        RECT 348.675 -10.365 349.005 -10.035 ;
        RECT 347.315 -10.365 347.645 -10.035 ;
        RECT 345.955 -10.365 346.285 -10.035 ;
        RECT 344.595 -10.365 344.925 -10.035 ;
        RECT 343.235 -10.365 343.565 -10.035 ;
        RECT 341.875 -10.365 342.205 -10.035 ;
        RECT 340.515 -10.365 340.845 -10.035 ;
        RECT 339.155 -10.365 339.485 -10.035 ;
        RECT 337.795 -10.365 338.125 -10.035 ;
        RECT 336.435 -10.365 336.765 -10.035 ;
        RECT 335.075 -10.365 335.405 -10.035 ;
        RECT 333.715 -10.365 334.045 -10.035 ;
        RECT 332.355 -10.365 332.685 -10.035 ;
        RECT 330.995 -10.365 331.325 -10.035 ;
        RECT 329.635 -10.365 329.965 -10.035 ;
        RECT 328.275 -10.365 328.605 -10.035 ;
        RECT 326.915 -10.365 327.245 -10.035 ;
        RECT 325.555 -10.365 325.885 -10.035 ;
        RECT 324.195 -10.365 324.525 -10.035 ;
        RECT 322.835 -10.365 323.165 -10.035 ;
        RECT 321.475 -10.365 321.805 -10.035 ;
        RECT 320.115 -10.365 320.445 -10.035 ;
        RECT 318.755 -10.365 319.085 -10.035 ;
        RECT 317.395 -10.365 317.725 -10.035 ;
        RECT 316.035 -10.365 316.365 -10.035 ;
        RECT 314.675 -10.365 315.005 -10.035 ;
        RECT 313.315 -10.365 313.645 -10.035 ;
        RECT 311.955 -10.365 312.285 -10.035 ;
        RECT 310.595 -10.365 310.925 -10.035 ;
        RECT 309.235 -10.365 309.565 -10.035 ;
        RECT 307.875 -10.365 308.205 -10.035 ;
        RECT 306.515 -10.365 306.845 -10.035 ;
        RECT 305.155 -10.365 305.485 -10.035 ;
        RECT 303.795 -10.365 304.125 -10.035 ;
        RECT 302.435 -10.365 302.765 -10.035 ;
        RECT 301.075 -10.365 301.405 -10.035 ;
        RECT 299.715 -10.365 300.045 -10.035 ;
        RECT 298.355 -10.365 298.685 -10.035 ;
        RECT 296.995 -10.365 297.325 -10.035 ;
        RECT 295.635 -10.365 295.965 -10.035 ;
        RECT 294.275 -10.365 294.605 -10.035 ;
        RECT 292.915 -10.365 293.245 -10.035 ;
        RECT 291.555 -10.365 291.885 -10.035 ;
        RECT 290.195 -10.365 290.525 -10.035 ;
        RECT 288.835 -10.365 289.165 -10.035 ;
        RECT 287.475 -10.365 287.805 -10.035 ;
        RECT 286.115 -10.365 286.445 -10.035 ;
        RECT 284.755 -10.365 285.085 -10.035 ;
        RECT 283.395 -10.365 283.725 -10.035 ;
        RECT 282.035 -10.365 282.365 -10.035 ;
        RECT 280.675 -10.365 281.005 -10.035 ;
        RECT 279.315 -10.365 279.645 -10.035 ;
        RECT 277.955 -10.365 278.285 -10.035 ;
        RECT 276.595 -10.365 276.925 -10.035 ;
        RECT 275.235 -10.365 275.565 -10.035 ;
        RECT 273.875 -10.365 274.205 -10.035 ;
        RECT 272.515 -10.365 272.845 -10.035 ;
        RECT 271.155 -10.365 271.485 -10.035 ;
        RECT 269.795 -10.365 270.125 -10.035 ;
        RECT 268.435 -10.365 268.765 -10.035 ;
        RECT 267.075 -10.365 267.405 -10.035 ;
        RECT 265.715 -10.365 266.045 -10.035 ;
        RECT 264.355 -10.365 264.685 -10.035 ;
        RECT 262.995 -10.365 263.325 -10.035 ;
        RECT 261.635 -10.365 261.965 -10.035 ;
        RECT 260.275 -10.365 260.605 -10.035 ;
        RECT 258.915 -10.365 259.245 -10.035 ;
        RECT 257.555 -10.365 257.885 -10.035 ;
        RECT 256.195 -10.365 256.525 -10.035 ;
        RECT 254.835 -10.365 255.165 -10.035 ;
        RECT 253.475 -10.365 253.805 -10.035 ;
        RECT 252.115 -10.365 252.445 -10.035 ;
        RECT 250.755 -10.365 251.085 -10.035 ;
        RECT 249.395 -10.365 249.725 -10.035 ;
        RECT 248.035 -10.365 248.365 -10.035 ;
        RECT 246.675 -10.365 247.005 -10.035 ;
        RECT 245.315 -10.365 245.645 -10.035 ;
        RECT 243.955 -10.365 244.285 -10.035 ;
        RECT 242.595 -10.365 242.925 -10.035 ;
        RECT 241.235 -10.365 241.565 -10.035 ;
        RECT 239.875 -10.365 240.205 -10.035 ;
        RECT 238.515 -10.365 238.845 -10.035 ;
        RECT 237.155 -10.365 237.485 -10.035 ;
        RECT 235.795 -10.365 236.125 -10.035 ;
        RECT 234.435 -10.365 234.765 -10.035 ;
        RECT 233.075 -10.365 233.405 -10.035 ;
        RECT 231.715 -10.365 232.045 -10.035 ;
        RECT 230.355 -10.365 230.685 -10.035 ;
        RECT 228.995 -10.365 229.325 -10.035 ;
        RECT 227.635 -10.365 227.965 -10.035 ;
        RECT 226.275 -10.365 226.605 -10.035 ;
        RECT 224.915 -10.365 225.245 -10.035 ;
        RECT 223.555 -10.365 223.885 -10.035 ;
        RECT 222.195 -10.365 222.525 -10.035 ;
        RECT 220.835 -10.365 221.165 -10.035 ;
        RECT 219.475 -10.365 219.805 -10.035 ;
        RECT 218.115 -10.365 218.445 -10.035 ;
        RECT 216.755 -10.365 217.085 -10.035 ;
        RECT 215.395 -10.365 215.725 -10.035 ;
        RECT 214.035 -10.365 214.365 -10.035 ;
        RECT 212.675 -10.365 213.005 -10.035 ;
        RECT 211.315 -10.365 211.645 -10.035 ;
        RECT 209.955 -10.365 210.285 -10.035 ;
        RECT 208.595 -10.365 208.925 -10.035 ;
        RECT 207.235 -10.365 207.565 -10.035 ;
        RECT 205.875 -10.365 206.205 -10.035 ;
        RECT 204.515 -10.365 204.845 -10.035 ;
        RECT 203.155 -10.365 203.485 -10.035 ;
        RECT 201.795 -10.365 202.125 -10.035 ;
        RECT 200.435 -10.365 200.765 -10.035 ;
        RECT 199.075 -10.365 199.405 -10.035 ;
        RECT 197.715 -10.365 198.045 -10.035 ;
        RECT 196.355 -10.365 196.685 -10.035 ;
        RECT 194.995 -10.365 195.325 -10.035 ;
        RECT 193.635 -10.365 193.965 -10.035 ;
        RECT 192.275 -10.365 192.605 -10.035 ;
        RECT 190.915 -10.365 191.245 -10.035 ;
        RECT 189.555 -10.365 189.885 -10.035 ;
        RECT 188.195 -10.365 188.525 -10.035 ;
        RECT 186.835 -10.365 187.165 -10.035 ;
        RECT 185.475 -10.365 185.805 -10.035 ;
        RECT 184.115 -10.365 184.445 -10.035 ;
        RECT 182.755 -10.365 183.085 -10.035 ;
        RECT 181.395 -10.365 181.725 -10.035 ;
        RECT 180.035 -10.365 180.365 -10.035 ;
        RECT 178.675 -10.365 179.005 -10.035 ;
        RECT 177.315 -10.365 177.645 -10.035 ;
        RECT 175.955 -10.365 176.285 -10.035 ;
        RECT 174.595 -10.365 174.925 -10.035 ;
        RECT 173.235 -10.365 173.565 -10.035 ;
        RECT 171.875 -10.365 172.205 -10.035 ;
        RECT 170.515 -10.365 170.845 -10.035 ;
        RECT 169.155 -10.365 169.485 -10.035 ;
        RECT 167.795 -10.365 168.125 -10.035 ;
        RECT 166.435 -10.365 166.765 -10.035 ;
        RECT 165.075 -10.365 165.405 -10.035 ;
        RECT 163.715 -10.365 164.045 -10.035 ;
        RECT 162.355 -10.365 162.685 -10.035 ;
        RECT 160.995 -10.365 161.325 -10.035 ;
        RECT 159.635 -10.365 159.965 -10.035 ;
        RECT 158.275 -10.365 158.605 -10.035 ;
        RECT 156.915 -10.365 157.245 -10.035 ;
        RECT 155.555 -10.365 155.885 -10.035 ;
        RECT 154.195 -10.365 154.525 -10.035 ;
        RECT 152.835 -10.365 153.165 -10.035 ;
        RECT 151.475 -10.365 151.805 -10.035 ;
        RECT 150.115 -10.365 150.445 -10.035 ;
        RECT 148.755 -10.365 149.085 -10.035 ;
        RECT 147.395 -10.365 147.725 -10.035 ;
        RECT 146.035 -10.365 146.365 -10.035 ;
        RECT 144.675 -10.365 145.005 -10.035 ;
        RECT 143.315 -10.365 143.645 -10.035 ;
        RECT 141.955 -10.365 142.285 -10.035 ;
        RECT 140.595 -10.365 140.925 -10.035 ;
        RECT 139.235 -10.365 139.565 -10.035 ;
        RECT 137.875 -10.365 138.205 -10.035 ;
        RECT 136.515 -10.365 136.845 -10.035 ;
        RECT 135.155 -10.365 135.485 -10.035 ;
        RECT 133.795 -10.365 134.125 -10.035 ;
        RECT 132.435 -10.365 132.765 -10.035 ;
        RECT 131.075 -10.365 131.405 -10.035 ;
        RECT 129.715 -10.365 130.045 -10.035 ;
        RECT 128.355 -10.365 128.685 -10.035 ;
        RECT 126.995 -10.365 127.325 -10.035 ;
        RECT 125.635 -10.365 125.965 -10.035 ;
        RECT 124.275 -10.365 124.605 -10.035 ;
        RECT 122.915 -10.365 123.245 -10.035 ;
        RECT 121.555 -10.365 121.885 -10.035 ;
        RECT 120.195 -10.365 120.525 -10.035 ;
        RECT 118.835 -10.365 119.165 -10.035 ;
        RECT 117.475 -10.365 117.805 -10.035 ;
        RECT 116.115 -10.365 116.445 -10.035 ;
        RECT 114.755 -10.365 115.085 -10.035 ;
        RECT 113.395 -10.365 113.725 -10.035 ;
        RECT 112.035 -10.365 112.365 -10.035 ;
        RECT 110.675 -10.365 111.005 -10.035 ;
        RECT 109.315 -10.365 109.645 -10.035 ;
        RECT 107.955 -10.365 108.285 -10.035 ;
        RECT 106.595 -10.365 106.925 -10.035 ;
        RECT 105.235 -10.365 105.565 -10.035 ;
        RECT 103.875 -10.365 104.205 -10.035 ;
        RECT 102.515 -10.365 102.845 -10.035 ;
        RECT 101.155 -10.365 101.485 -10.035 ;
        RECT 99.795 -10.365 100.125 -10.035 ;
        RECT 98.435 -10.365 98.765 -10.035 ;
        RECT 97.075 -10.365 97.405 -10.035 ;
        RECT 95.715 -10.365 96.045 -10.035 ;
        RECT 94.355 -10.365 94.685 -10.035 ;
        RECT 92.995 -10.365 93.325 -10.035 ;
        RECT 91.635 -10.365 91.965 -10.035 ;
        RECT 90.275 -10.365 90.605 -10.035 ;
        RECT 88.915 -10.365 89.245 -10.035 ;
        RECT 87.555 -10.365 87.885 -10.035 ;
        RECT 86.195 -10.365 86.525 -10.035 ;
        RECT 84.835 -10.365 85.165 -10.035 ;
        RECT 83.475 -10.365 83.805 -10.035 ;
        RECT 82.115 -10.365 82.445 -10.035 ;
        RECT 80.755 -10.365 81.085 -10.035 ;
        RECT 79.395 -10.365 79.725 -10.035 ;
        RECT 78.035 -10.365 78.365 -10.035 ;
        RECT 76.675 -10.365 77.005 -10.035 ;
        RECT 75.315 -10.365 75.645 -10.035 ;
        RECT 73.955 -10.365 74.285 -10.035 ;
        RECT 72.595 -10.365 72.925 -10.035 ;
        RECT 71.235 -10.365 71.565 -10.035 ;
        RECT 69.875 -10.365 70.205 -10.035 ;
        RECT 68.515 -10.365 68.845 -10.035 ;
        RECT 67.155 -10.365 67.485 -10.035 ;
        RECT 65.795 -10.365 66.125 -10.035 ;
        RECT 64.435 -10.365 64.765 -10.035 ;
        RECT 63.075 -10.365 63.405 -10.035 ;
        RECT 61.715 -10.365 62.045 -10.035 ;
        RECT 60.355 -10.365 60.685 -10.035 ;
        RECT 58.995 -10.365 59.325 -10.035 ;
        RECT 57.635 -10.365 57.965 -10.035 ;
        RECT 56.275 -10.365 56.605 -10.035 ;
        RECT 54.915 -10.365 55.245 -10.035 ;
        RECT 53.555 -10.365 53.885 -10.035 ;
        RECT 52.195 -10.365 52.525 -10.035 ;
        RECT 50.835 -10.365 51.165 -10.035 ;
        RECT 49.475 -10.365 49.805 -10.035 ;
        RECT 48.115 -10.365 48.445 -10.035 ;
        RECT 46.755 -10.365 47.085 -10.035 ;
        RECT 45.395 -10.365 45.725 -10.035 ;
        RECT 44.035 -10.365 44.365 -10.035 ;
        RECT 42.675 -10.365 43.005 -10.035 ;
        RECT 41.315 -10.365 41.645 -10.035 ;
        RECT 39.955 -10.365 40.285 -10.035 ;
        RECT 38.595 -10.365 38.925 -10.035 ;
        RECT 37.235 -10.365 37.565 -10.035 ;
        RECT 35.875 -10.365 36.205 -10.035 ;
        RECT 34.515 -10.365 34.845 -10.035 ;
        RECT 33.155 -10.365 33.485 -10.035 ;
        RECT 31.795 -10.365 32.125 -10.035 ;
        RECT 30.435 -10.365 30.765 -10.035 ;
        RECT 29.075 -10.365 29.405 -10.035 ;
        RECT 27.715 -10.365 28.045 -10.035 ;
        RECT 26.355 -10.365 26.685 -10.035 ;
        RECT 24.995 -10.365 25.325 -10.035 ;
        RECT 23.635 -10.365 23.965 -10.035 ;
        RECT 22.275 -10.365 22.605 -10.035 ;
        RECT 20.915 -10.365 21.245 -10.035 ;
        RECT 19.555 -10.365 19.885 -10.035 ;
        RECT 18.195 -10.365 18.525 -10.035 ;
        RECT 16.835 -10.365 17.165 -10.035 ;
        RECT 15.475 -10.365 15.805 -10.035 ;
        RECT 14.115 -10.365 14.445 -10.035 ;
        RECT 12.755 -10.365 13.085 -10.035 ;
        RECT 11.395 -10.365 11.725 -10.035 ;
        RECT 10.035 -10.365 10.365 -10.035 ;
        RECT 8.675 -10.365 9.005 -10.035 ;
        RECT 7.315 -10.365 7.645 -10.035 ;
        RECT 5.955 -10.365 6.285 -10.035 ;
        RECT 4.595 -10.365 4.925 -10.035 ;
        RECT 3.235 -10.365 3.565 -10.035 ;
        RECT 1.875 -10.365 2.205 -10.035 ;
        RECT 0.515 -10.365 0.845 -10.035 ;
        RECT -0.845 -10.365 -0.515 -10.035 ;
        RECT 678.125 -10.36 954.88 -10.04 ;
        RECT 953.875 -10.365 954.205 -10.035 ;
        RECT 952.515 -10.365 952.845 -10.035 ;
        RECT 951.155 -10.365 951.485 -10.035 ;
        RECT 949.795 -10.365 950.125 -10.035 ;
        RECT 948.435 -10.365 948.765 -10.035 ;
        RECT 947.075 -10.365 947.405 -10.035 ;
        RECT 945.715 -10.365 946.045 -10.035 ;
        RECT 944.355 -10.365 944.685 -10.035 ;
        RECT 942.995 -10.365 943.325 -10.035 ;
        RECT 941.635 -10.365 941.965 -10.035 ;
        RECT 940.275 -10.365 940.605 -10.035 ;
        RECT 938.915 -10.365 939.245 -10.035 ;
        RECT 937.555 -10.365 937.885 -10.035 ;
        RECT 936.195 -10.365 936.525 -10.035 ;
        RECT 934.835 -10.365 935.165 -10.035 ;
        RECT 933.475 -10.365 933.805 -10.035 ;
        RECT 932.115 -10.365 932.445 -10.035 ;
        RECT 930.755 -10.365 931.085 -10.035 ;
        RECT 929.395 -10.365 929.725 -10.035 ;
        RECT 928.035 -10.365 928.365 -10.035 ;
        RECT 926.675 -10.365 927.005 -10.035 ;
        RECT 925.315 -10.365 925.645 -10.035 ;
        RECT 923.955 -10.365 924.285 -10.035 ;
        RECT 922.595 -10.365 922.925 -10.035 ;
        RECT 921.235 -10.365 921.565 -10.035 ;
        RECT 919.875 -10.365 920.205 -10.035 ;
        RECT 918.515 -10.365 918.845 -10.035 ;
        RECT 917.155 -10.365 917.485 -10.035 ;
        RECT 915.795 -10.365 916.125 -10.035 ;
        RECT 914.435 -10.365 914.765 -10.035 ;
        RECT 913.075 -10.365 913.405 -10.035 ;
        RECT 911.715 -10.365 912.045 -10.035 ;
        RECT 910.355 -10.365 910.685 -10.035 ;
        RECT 908.995 -10.365 909.325 -10.035 ;
        RECT 907.635 -10.365 907.965 -10.035 ;
        RECT 906.275 -10.365 906.605 -10.035 ;
        RECT 904.915 -10.365 905.245 -10.035 ;
        RECT 903.555 -10.365 903.885 -10.035 ;
        RECT 902.195 -10.365 902.525 -10.035 ;
        RECT 900.835 -10.365 901.165 -10.035 ;
        RECT 899.475 -10.365 899.805 -10.035 ;
        RECT 898.115 -10.365 898.445 -10.035 ;
        RECT 896.755 -10.365 897.085 -10.035 ;
        RECT 895.395 -10.365 895.725 -10.035 ;
        RECT 894.035 -10.365 894.365 -10.035 ;
        RECT 892.675 -10.365 893.005 -10.035 ;
        RECT 891.315 -10.365 891.645 -10.035 ;
        RECT 889.955 -10.365 890.285 -10.035 ;
        RECT 888.595 -10.365 888.925 -10.035 ;
        RECT 887.235 -10.365 887.565 -10.035 ;
        RECT 885.875 -10.365 886.205 -10.035 ;
        RECT 884.515 -10.365 884.845 -10.035 ;
        RECT 883.155 -10.365 883.485 -10.035 ;
        RECT 881.795 -10.365 882.125 -10.035 ;
        RECT 880.435 -10.365 880.765 -10.035 ;
        RECT 879.075 -10.365 879.405 -10.035 ;
        RECT 877.715 -10.365 878.045 -10.035 ;
        RECT 876.355 -10.365 876.685 -10.035 ;
        RECT 874.995 -10.365 875.325 -10.035 ;
        RECT 873.635 -10.365 873.965 -10.035 ;
        RECT 872.275 -10.365 872.605 -10.035 ;
        RECT 870.915 -10.365 871.245 -10.035 ;
        RECT 869.555 -10.365 869.885 -10.035 ;
        RECT 868.195 -10.365 868.525 -10.035 ;
        RECT 866.835 -10.365 867.165 -10.035 ;
        RECT 865.475 -10.365 865.805 -10.035 ;
        RECT 864.115 -10.365 864.445 -10.035 ;
        RECT 862.755 -10.365 863.085 -10.035 ;
        RECT 861.395 -10.365 861.725 -10.035 ;
        RECT 860.035 -10.365 860.365 -10.035 ;
        RECT 858.675 -10.365 859.005 -10.035 ;
        RECT 857.315 -10.365 857.645 -10.035 ;
        RECT 855.955 -10.365 856.285 -10.035 ;
        RECT 854.595 -10.365 854.925 -10.035 ;
        RECT 853.235 -10.365 853.565 -10.035 ;
        RECT 851.875 -10.365 852.205 -10.035 ;
        RECT 850.515 -10.365 850.845 -10.035 ;
        RECT 849.155 -10.365 849.485 -10.035 ;
        RECT 847.795 -10.365 848.125 -10.035 ;
        RECT 846.435 -10.365 846.765 -10.035 ;
        RECT 845.075 -10.365 845.405 -10.035 ;
        RECT 843.715 -10.365 844.045 -10.035 ;
        RECT 842.355 -10.365 842.685 -10.035 ;
        RECT 840.995 -10.365 841.325 -10.035 ;
        RECT 839.635 -10.365 839.965 -10.035 ;
        RECT 838.275 -10.365 838.605 -10.035 ;
        RECT 836.915 -10.365 837.245 -10.035 ;
        RECT 835.555 -10.365 835.885 -10.035 ;
        RECT 834.195 -10.365 834.525 -10.035 ;
        RECT 832.835 -10.365 833.165 -10.035 ;
        RECT 831.475 -10.365 831.805 -10.035 ;
        RECT 830.115 -10.365 830.445 -10.035 ;
        RECT 828.755 -10.365 829.085 -10.035 ;
        RECT 827.395 -10.365 827.725 -10.035 ;
        RECT 826.035 -10.365 826.365 -10.035 ;
        RECT 824.675 -10.365 825.005 -10.035 ;
        RECT 823.315 -10.365 823.645 -10.035 ;
        RECT 821.955 -10.365 822.285 -10.035 ;
        RECT 820.595 -10.365 820.925 -10.035 ;
        RECT 819.235 -10.365 819.565 -10.035 ;
        RECT 817.875 -10.365 818.205 -10.035 ;
        RECT 816.515 -10.365 816.845 -10.035 ;
        RECT 815.155 -10.365 815.485 -10.035 ;
        RECT 813.795 -10.365 814.125 -10.035 ;
        RECT 812.435 -10.365 812.765 -10.035 ;
        RECT 811.075 -10.365 811.405 -10.035 ;
        RECT 809.715 -10.365 810.045 -10.035 ;
        RECT 808.355 -10.365 808.685 -10.035 ;
        RECT 806.995 -10.365 807.325 -10.035 ;
        RECT 805.635 -10.365 805.965 -10.035 ;
        RECT 804.275 -10.365 804.605 -10.035 ;
        RECT 802.915 -10.365 803.245 -10.035 ;
        RECT 801.555 -10.365 801.885 -10.035 ;
        RECT 800.195 -10.365 800.525 -10.035 ;
        RECT 798.835 -10.365 799.165 -10.035 ;
        RECT 797.475 -10.365 797.805 -10.035 ;
        RECT 796.115 -10.365 796.445 -10.035 ;
        RECT 794.755 -10.365 795.085 -10.035 ;
        RECT 793.395 -10.365 793.725 -10.035 ;
        RECT 792.035 -10.365 792.365 -10.035 ;
        RECT 790.675 -10.365 791.005 -10.035 ;
        RECT 789.315 -10.365 789.645 -10.035 ;
        RECT 787.955 -10.365 788.285 -10.035 ;
        RECT 786.595 -10.365 786.925 -10.035 ;
        RECT 785.235 -10.365 785.565 -10.035 ;
        RECT 783.875 -10.365 784.205 -10.035 ;
        RECT 782.515 -10.365 782.845 -10.035 ;
        RECT 781.155 -10.365 781.485 -10.035 ;
        RECT 779.795 -10.365 780.125 -10.035 ;
        RECT 778.435 -10.365 778.765 -10.035 ;
        RECT 777.075 -10.365 777.405 -10.035 ;
        RECT 775.715 -10.365 776.045 -10.035 ;
        RECT 774.355 -10.365 774.685 -10.035 ;
        RECT 772.995 -10.365 773.325 -10.035 ;
        RECT 771.635 -10.365 771.965 -10.035 ;
        RECT 770.275 -10.365 770.605 -10.035 ;
        RECT 768.915 -10.365 769.245 -10.035 ;
        RECT 767.555 -10.365 767.885 -10.035 ;
        RECT 766.195 -10.365 766.525 -10.035 ;
        RECT 764.835 -10.365 765.165 -10.035 ;
        RECT 763.475 -10.365 763.805 -10.035 ;
        RECT 762.115 -10.365 762.445 -10.035 ;
        RECT 760.755 -10.365 761.085 -10.035 ;
        RECT 759.395 -10.365 759.725 -10.035 ;
        RECT 758.035 -10.365 758.365 -10.035 ;
        RECT 756.675 -10.365 757.005 -10.035 ;
        RECT 755.315 -10.365 755.645 -10.035 ;
        RECT 753.955 -10.365 754.285 -10.035 ;
        RECT 752.595 -10.365 752.925 -10.035 ;
        RECT 751.235 -10.365 751.565 -10.035 ;
        RECT 749.875 -10.365 750.205 -10.035 ;
        RECT 748.515 -10.365 748.845 -10.035 ;
        RECT 747.155 -10.365 747.485 -10.035 ;
        RECT 745.795 -10.365 746.125 -10.035 ;
        RECT 744.435 -10.365 744.765 -10.035 ;
        RECT 743.075 -10.365 743.405 -10.035 ;
        RECT 741.715 -10.365 742.045 -10.035 ;
        RECT 740.355 -10.365 740.685 -10.035 ;
        RECT 738.995 -10.365 739.325 -10.035 ;
        RECT 737.635 -10.365 737.965 -10.035 ;
        RECT 736.275 -10.365 736.605 -10.035 ;
        RECT 734.915 -10.365 735.245 -10.035 ;
        RECT 733.555 -10.365 733.885 -10.035 ;
        RECT 732.195 -10.365 732.525 -10.035 ;
        RECT 730.835 -10.365 731.165 -10.035 ;
        RECT 729.475 -10.365 729.805 -10.035 ;
        RECT 728.115 -10.365 728.445 -10.035 ;
        RECT 726.755 -10.365 727.085 -10.035 ;
        RECT 725.395 -10.365 725.725 -10.035 ;
        RECT 724.035 -10.365 724.365 -10.035 ;
        RECT 722.675 -10.365 723.005 -10.035 ;
        RECT 721.315 -10.365 721.645 -10.035 ;
        RECT 719.955 -10.365 720.285 -10.035 ;
        RECT 718.595 -10.365 718.925 -10.035 ;
        RECT 717.235 -10.365 717.565 -10.035 ;
        RECT 715.875 -10.365 716.205 -10.035 ;
        RECT 714.515 -10.365 714.845 -10.035 ;
        RECT 713.155 -10.365 713.485 -10.035 ;
        RECT 711.795 -10.365 712.125 -10.035 ;
        RECT 710.435 -10.365 710.765 -10.035 ;
        RECT 709.075 -10.365 709.405 -10.035 ;
        RECT 707.715 -10.365 708.045 -10.035 ;
        RECT 706.355 -10.365 706.685 -10.035 ;
        RECT 704.995 -10.365 705.325 -10.035 ;
        RECT 703.635 -10.365 703.965 -10.035 ;
        RECT 702.275 -10.365 702.605 -10.035 ;
        RECT 700.915 -10.365 701.245 -10.035 ;
        RECT 699.555 -10.365 699.885 -10.035 ;
        RECT 698.195 -10.365 698.525 -10.035 ;
        RECT 696.835 -10.365 697.165 -10.035 ;
        RECT 695.475 -10.365 695.805 -10.035 ;
        RECT 694.115 -10.365 694.445 -10.035 ;
        RECT 692.755 -10.365 693.085 -10.035 ;
        RECT 691.395 -10.365 691.725 -10.035 ;
        RECT 690.035 -10.365 690.365 -10.035 ;
        RECT 688.675 -10.365 689.005 -10.035 ;
        RECT 687.315 -10.365 687.645 -10.035 ;
        RECT 685.955 -10.365 686.285 -10.035 ;
        RECT 684.595 -10.365 684.925 -10.035 ;
        RECT 683.235 -10.365 683.565 -10.035 ;
        RECT 681.875 -10.365 682.205 -10.035 ;
        RECT 680.515 -10.365 680.845 -10.035 ;
        RECT 679.155 -10.365 679.485 -10.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -11.725 128.685 -11.395 ;
        RECT 126.995 -11.725 127.325 -11.395 ;
        RECT 125.635 -11.725 125.965 -11.395 ;
        RECT 124.275 -11.725 124.605 -11.395 ;
        RECT 122.915 -11.725 123.245 -11.395 ;
        RECT 121.555 -11.725 121.885 -11.395 ;
        RECT 120.195 -11.725 120.525 -11.395 ;
        RECT 118.835 -11.725 119.165 -11.395 ;
        RECT 117.475 -11.725 117.805 -11.395 ;
        RECT 116.115 -11.725 116.445 -11.395 ;
        RECT 114.755 -11.725 115.085 -11.395 ;
        RECT 113.395 -11.725 113.725 -11.395 ;
        RECT 112.035 -11.725 112.365 -11.395 ;
        RECT 110.675 -11.725 111.005 -11.395 ;
        RECT 109.315 -11.725 109.645 -11.395 ;
        RECT 107.955 -11.725 108.285 -11.395 ;
        RECT 106.595 -11.725 106.925 -11.395 ;
        RECT 105.235 -11.725 105.565 -11.395 ;
        RECT 103.875 -11.725 104.205 -11.395 ;
        RECT 102.515 -11.725 102.845 -11.395 ;
        RECT 101.155 -11.725 101.485 -11.395 ;
        RECT 99.795 -11.725 100.125 -11.395 ;
        RECT 98.435 -11.725 98.765 -11.395 ;
        RECT 97.075 -11.725 97.405 -11.395 ;
        RECT 95.715 -11.725 96.045 -11.395 ;
        RECT 94.355 -11.725 94.685 -11.395 ;
        RECT 92.995 -11.725 93.325 -11.395 ;
        RECT 91.635 -11.725 91.965 -11.395 ;
        RECT 90.275 -11.725 90.605 -11.395 ;
        RECT 88.915 -11.725 89.245 -11.395 ;
        RECT 87.555 -11.725 87.885 -11.395 ;
        RECT 86.195 -11.725 86.525 -11.395 ;
        RECT 84.835 -11.725 85.165 -11.395 ;
        RECT 83.475 -11.725 83.805 -11.395 ;
        RECT 82.115 -11.725 82.445 -11.395 ;
        RECT 80.755 -11.725 81.085 -11.395 ;
        RECT 79.395 -11.725 79.725 -11.395 ;
        RECT 78.035 -11.725 78.365 -11.395 ;
        RECT 76.675 -11.725 77.005 -11.395 ;
        RECT 75.315 -11.725 75.645 -11.395 ;
        RECT 73.955 -11.725 74.285 -11.395 ;
        RECT 72.595 -11.725 72.925 -11.395 ;
        RECT 71.235 -11.725 71.565 -11.395 ;
        RECT 69.875 -11.725 70.205 -11.395 ;
        RECT 68.515 -11.725 68.845 -11.395 ;
        RECT 67.155 -11.725 67.485 -11.395 ;
        RECT 65.795 -11.725 66.125 -11.395 ;
        RECT 64.435 -11.725 64.765 -11.395 ;
        RECT 63.075 -11.725 63.405 -11.395 ;
        RECT 61.715 -11.725 62.045 -11.395 ;
        RECT 60.355 -11.725 60.685 -11.395 ;
        RECT 58.995 -11.725 59.325 -11.395 ;
        RECT 57.635 -11.725 57.965 -11.395 ;
        RECT 56.275 -11.725 56.605 -11.395 ;
        RECT 54.915 -11.725 55.245 -11.395 ;
        RECT 53.555 -11.725 53.885 -11.395 ;
        RECT 52.195 -11.725 52.525 -11.395 ;
        RECT 50.835 -11.725 51.165 -11.395 ;
        RECT 49.475 -11.725 49.805 -11.395 ;
        RECT 48.115 -11.725 48.445 -11.395 ;
        RECT 46.755 -11.725 47.085 -11.395 ;
        RECT 45.395 -11.725 45.725 -11.395 ;
        RECT 44.035 -11.725 44.365 -11.395 ;
        RECT 42.675 -11.725 43.005 -11.395 ;
        RECT 41.315 -11.725 41.645 -11.395 ;
        RECT 39.955 -11.725 40.285 -11.395 ;
        RECT 38.595 -11.725 38.925 -11.395 ;
        RECT 37.235 -11.725 37.565 -11.395 ;
        RECT 35.875 -11.725 36.205 -11.395 ;
        RECT 34.515 -11.725 34.845 -11.395 ;
        RECT 33.155 -11.725 33.485 -11.395 ;
        RECT 31.795 -11.725 32.125 -11.395 ;
        RECT 30.435 -11.725 30.765 -11.395 ;
        RECT 29.075 -11.725 29.405 -11.395 ;
        RECT 27.715 -11.725 28.045 -11.395 ;
        RECT 26.355 -11.725 26.685 -11.395 ;
        RECT 24.995 -11.725 25.325 -11.395 ;
        RECT 23.635 -11.725 23.965 -11.395 ;
        RECT 22.275 -11.725 22.605 -11.395 ;
        RECT 20.915 -11.725 21.245 -11.395 ;
        RECT 19.555 -11.725 19.885 -11.395 ;
        RECT 18.195 -11.725 18.525 -11.395 ;
        RECT 16.835 -11.725 17.165 -11.395 ;
        RECT 15.475 -11.725 15.805 -11.395 ;
        RECT 14.115 -11.725 14.445 -11.395 ;
        RECT 12.755 -11.725 13.085 -11.395 ;
        RECT 11.395 -11.725 11.725 -11.395 ;
        RECT 10.035 -11.725 10.365 -11.395 ;
        RECT 8.675 -11.725 9.005 -11.395 ;
        RECT 7.315 -11.725 7.645 -11.395 ;
        RECT 5.955 -11.725 6.285 -11.395 ;
        RECT 4.595 -11.725 4.925 -11.395 ;
        RECT 3.235 -11.725 3.565 -11.395 ;
        RECT 1.875 -11.725 2.205 -11.395 ;
        RECT 0.515 -11.725 0.845 -11.395 ;
        RECT -0.845 -11.725 -0.515 -11.395 ;
        RECT 677.795 -11.725 678.125 -11.395 ;
        RECT -1.52 -11.72 678.125 -11.4 ;
        RECT 676.435 -11.725 676.765 -11.395 ;
        RECT 675.075 -11.725 675.405 -11.395 ;
        RECT 673.715 -11.725 674.045 -11.395 ;
        RECT 672.355 -11.725 672.685 -11.395 ;
        RECT 670.995 -11.725 671.325 -11.395 ;
        RECT 669.635 -11.725 669.965 -11.395 ;
        RECT 668.275 -11.725 668.605 -11.395 ;
        RECT 666.915 -11.725 667.245 -11.395 ;
        RECT 665.555 -11.725 665.885 -11.395 ;
        RECT 664.195 -11.725 664.525 -11.395 ;
        RECT 662.835 -11.725 663.165 -11.395 ;
        RECT 661.475 -11.725 661.805 -11.395 ;
        RECT 660.115 -11.725 660.445 -11.395 ;
        RECT 658.755 -11.725 659.085 -11.395 ;
        RECT 657.395 -11.725 657.725 -11.395 ;
        RECT 656.035 -11.725 656.365 -11.395 ;
        RECT 654.675 -11.725 655.005 -11.395 ;
        RECT 653.315 -11.725 653.645 -11.395 ;
        RECT 651.955 -11.725 652.285 -11.395 ;
        RECT 650.595 -11.725 650.925 -11.395 ;
        RECT 649.235 -11.725 649.565 -11.395 ;
        RECT 647.875 -11.725 648.205 -11.395 ;
        RECT 646.515 -11.725 646.845 -11.395 ;
        RECT 645.155 -11.725 645.485 -11.395 ;
        RECT 643.795 -11.725 644.125 -11.395 ;
        RECT 642.435 -11.725 642.765 -11.395 ;
        RECT 641.075 -11.725 641.405 -11.395 ;
        RECT 639.715 -11.725 640.045 -11.395 ;
        RECT 638.355 -11.725 638.685 -11.395 ;
        RECT 636.995 -11.725 637.325 -11.395 ;
        RECT 635.635 -11.725 635.965 -11.395 ;
        RECT 634.275 -11.725 634.605 -11.395 ;
        RECT 632.915 -11.725 633.245 -11.395 ;
        RECT 631.555 -11.725 631.885 -11.395 ;
        RECT 630.195 -11.725 630.525 -11.395 ;
        RECT 628.835 -11.725 629.165 -11.395 ;
        RECT 627.475 -11.725 627.805 -11.395 ;
        RECT 626.115 -11.725 626.445 -11.395 ;
        RECT 624.755 -11.725 625.085 -11.395 ;
        RECT 623.395 -11.725 623.725 -11.395 ;
        RECT 622.035 -11.725 622.365 -11.395 ;
        RECT 620.675 -11.725 621.005 -11.395 ;
        RECT 619.315 -11.725 619.645 -11.395 ;
        RECT 617.955 -11.725 618.285 -11.395 ;
        RECT 616.595 -11.725 616.925 -11.395 ;
        RECT 615.235 -11.725 615.565 -11.395 ;
        RECT 613.875 -11.725 614.205 -11.395 ;
        RECT 612.515 -11.725 612.845 -11.395 ;
        RECT 611.155 -11.725 611.485 -11.395 ;
        RECT 609.795 -11.725 610.125 -11.395 ;
        RECT 608.435 -11.725 608.765 -11.395 ;
        RECT 607.075 -11.725 607.405 -11.395 ;
        RECT 605.715 -11.725 606.045 -11.395 ;
        RECT 604.355 -11.725 604.685 -11.395 ;
        RECT 602.995 -11.725 603.325 -11.395 ;
        RECT 601.635 -11.725 601.965 -11.395 ;
        RECT 600.275 -11.725 600.605 -11.395 ;
        RECT 598.915 -11.725 599.245 -11.395 ;
        RECT 597.555 -11.725 597.885 -11.395 ;
        RECT 596.195 -11.725 596.525 -11.395 ;
        RECT 594.835 -11.725 595.165 -11.395 ;
        RECT 593.475 -11.725 593.805 -11.395 ;
        RECT 592.115 -11.725 592.445 -11.395 ;
        RECT 590.755 -11.725 591.085 -11.395 ;
        RECT 589.395 -11.725 589.725 -11.395 ;
        RECT 588.035 -11.725 588.365 -11.395 ;
        RECT 586.675 -11.725 587.005 -11.395 ;
        RECT 585.315 -11.725 585.645 -11.395 ;
        RECT 583.955 -11.725 584.285 -11.395 ;
        RECT 582.595 -11.725 582.925 -11.395 ;
        RECT 581.235 -11.725 581.565 -11.395 ;
        RECT 579.875 -11.725 580.205 -11.395 ;
        RECT 578.515 -11.725 578.845 -11.395 ;
        RECT 577.155 -11.725 577.485 -11.395 ;
        RECT 575.795 -11.725 576.125 -11.395 ;
        RECT 574.435 -11.725 574.765 -11.395 ;
        RECT 573.075 -11.725 573.405 -11.395 ;
        RECT 571.715 -11.725 572.045 -11.395 ;
        RECT 570.355 -11.725 570.685 -11.395 ;
        RECT 568.995 -11.725 569.325 -11.395 ;
        RECT 567.635 -11.725 567.965 -11.395 ;
        RECT 566.275 -11.725 566.605 -11.395 ;
        RECT 564.915 -11.725 565.245 -11.395 ;
        RECT 563.555 -11.725 563.885 -11.395 ;
        RECT 562.195 -11.725 562.525 -11.395 ;
        RECT 560.835 -11.725 561.165 -11.395 ;
        RECT 559.475 -11.725 559.805 -11.395 ;
        RECT 558.115 -11.725 558.445 -11.395 ;
        RECT 556.755 -11.725 557.085 -11.395 ;
        RECT 555.395 -11.725 555.725 -11.395 ;
        RECT 554.035 -11.725 554.365 -11.395 ;
        RECT 552.675 -11.725 553.005 -11.395 ;
        RECT 551.315 -11.725 551.645 -11.395 ;
        RECT 549.955 -11.725 550.285 -11.395 ;
        RECT 548.595 -11.725 548.925 -11.395 ;
        RECT 547.235 -11.725 547.565 -11.395 ;
        RECT 545.875 -11.725 546.205 -11.395 ;
        RECT 544.515 -11.725 544.845 -11.395 ;
        RECT 543.155 -11.725 543.485 -11.395 ;
        RECT 541.795 -11.725 542.125 -11.395 ;
        RECT 540.435 -11.725 540.765 -11.395 ;
        RECT 539.075 -11.725 539.405 -11.395 ;
        RECT 537.715 -11.725 538.045 -11.395 ;
        RECT 536.355 -11.725 536.685 -11.395 ;
        RECT 534.995 -11.725 535.325 -11.395 ;
        RECT 533.635 -11.725 533.965 -11.395 ;
        RECT 532.275 -11.725 532.605 -11.395 ;
        RECT 530.915 -11.725 531.245 -11.395 ;
        RECT 529.555 -11.725 529.885 -11.395 ;
        RECT 528.195 -11.725 528.525 -11.395 ;
        RECT 526.835 -11.725 527.165 -11.395 ;
        RECT 525.475 -11.725 525.805 -11.395 ;
        RECT 524.115 -11.725 524.445 -11.395 ;
        RECT 522.755 -11.725 523.085 -11.395 ;
        RECT 521.395 -11.725 521.725 -11.395 ;
        RECT 520.035 -11.725 520.365 -11.395 ;
        RECT 518.675 -11.725 519.005 -11.395 ;
        RECT 517.315 -11.725 517.645 -11.395 ;
        RECT 515.955 -11.725 516.285 -11.395 ;
        RECT 514.595 -11.725 514.925 -11.395 ;
        RECT 513.235 -11.725 513.565 -11.395 ;
        RECT 511.875 -11.725 512.205 -11.395 ;
        RECT 510.515 -11.725 510.845 -11.395 ;
        RECT 509.155 -11.725 509.485 -11.395 ;
        RECT 507.795 -11.725 508.125 -11.395 ;
        RECT 506.435 -11.725 506.765 -11.395 ;
        RECT 505.075 -11.725 505.405 -11.395 ;
        RECT 503.715 -11.725 504.045 -11.395 ;
        RECT 502.355 -11.725 502.685 -11.395 ;
        RECT 500.995 -11.725 501.325 -11.395 ;
        RECT 499.635 -11.725 499.965 -11.395 ;
        RECT 498.275 -11.725 498.605 -11.395 ;
        RECT 496.915 -11.725 497.245 -11.395 ;
        RECT 495.555 -11.725 495.885 -11.395 ;
        RECT 494.195 -11.725 494.525 -11.395 ;
        RECT 492.835 -11.725 493.165 -11.395 ;
        RECT 491.475 -11.725 491.805 -11.395 ;
        RECT 490.115 -11.725 490.445 -11.395 ;
        RECT 488.755 -11.725 489.085 -11.395 ;
        RECT 487.395 -11.725 487.725 -11.395 ;
        RECT 486.035 -11.725 486.365 -11.395 ;
        RECT 484.675 -11.725 485.005 -11.395 ;
        RECT 483.315 -11.725 483.645 -11.395 ;
        RECT 481.955 -11.725 482.285 -11.395 ;
        RECT 480.595 -11.725 480.925 -11.395 ;
        RECT 479.235 -11.725 479.565 -11.395 ;
        RECT 477.875 -11.725 478.205 -11.395 ;
        RECT 476.515 -11.725 476.845 -11.395 ;
        RECT 475.155 -11.725 475.485 -11.395 ;
        RECT 473.795 -11.725 474.125 -11.395 ;
        RECT 472.435 -11.725 472.765 -11.395 ;
        RECT 471.075 -11.725 471.405 -11.395 ;
        RECT 469.715 -11.725 470.045 -11.395 ;
        RECT 468.355 -11.725 468.685 -11.395 ;
        RECT 466.995 -11.725 467.325 -11.395 ;
        RECT 465.635 -11.725 465.965 -11.395 ;
        RECT 464.275 -11.725 464.605 -11.395 ;
        RECT 462.915 -11.725 463.245 -11.395 ;
        RECT 461.555 -11.725 461.885 -11.395 ;
        RECT 460.195 -11.725 460.525 -11.395 ;
        RECT 458.835 -11.725 459.165 -11.395 ;
        RECT 457.475 -11.725 457.805 -11.395 ;
        RECT 456.115 -11.725 456.445 -11.395 ;
        RECT 454.755 -11.725 455.085 -11.395 ;
        RECT 453.395 -11.725 453.725 -11.395 ;
        RECT 452.035 -11.725 452.365 -11.395 ;
        RECT 450.675 -11.725 451.005 -11.395 ;
        RECT 449.315 -11.725 449.645 -11.395 ;
        RECT 447.955 -11.725 448.285 -11.395 ;
        RECT 446.595 -11.725 446.925 -11.395 ;
        RECT 445.235 -11.725 445.565 -11.395 ;
        RECT 443.875 -11.725 444.205 -11.395 ;
        RECT 442.515 -11.725 442.845 -11.395 ;
        RECT 441.155 -11.725 441.485 -11.395 ;
        RECT 439.795 -11.725 440.125 -11.395 ;
        RECT 438.435 -11.725 438.765 -11.395 ;
        RECT 437.075 -11.725 437.405 -11.395 ;
        RECT 435.715 -11.725 436.045 -11.395 ;
        RECT 434.355 -11.725 434.685 -11.395 ;
        RECT 432.995 -11.725 433.325 -11.395 ;
        RECT 431.635 -11.725 431.965 -11.395 ;
        RECT 430.275 -11.725 430.605 -11.395 ;
        RECT 428.915 -11.725 429.245 -11.395 ;
        RECT 427.555 -11.725 427.885 -11.395 ;
        RECT 426.195 -11.725 426.525 -11.395 ;
        RECT 424.835 -11.725 425.165 -11.395 ;
        RECT 423.475 -11.725 423.805 -11.395 ;
        RECT 422.115 -11.725 422.445 -11.395 ;
        RECT 420.755 -11.725 421.085 -11.395 ;
        RECT 419.395 -11.725 419.725 -11.395 ;
        RECT 418.035 -11.725 418.365 -11.395 ;
        RECT 416.675 -11.725 417.005 -11.395 ;
        RECT 415.315 -11.725 415.645 -11.395 ;
        RECT 413.955 -11.725 414.285 -11.395 ;
        RECT 412.595 -11.725 412.925 -11.395 ;
        RECT 411.235 -11.725 411.565 -11.395 ;
        RECT 409.875 -11.725 410.205 -11.395 ;
        RECT 408.515 -11.725 408.845 -11.395 ;
        RECT 407.155 -11.725 407.485 -11.395 ;
        RECT 405.795 -11.725 406.125 -11.395 ;
        RECT 404.435 -11.725 404.765 -11.395 ;
        RECT 403.075 -11.725 403.405 -11.395 ;
        RECT 401.715 -11.725 402.045 -11.395 ;
        RECT 400.355 -11.725 400.685 -11.395 ;
        RECT 398.995 -11.725 399.325 -11.395 ;
        RECT 397.635 -11.725 397.965 -11.395 ;
        RECT 396.275 -11.725 396.605 -11.395 ;
        RECT 394.915 -11.725 395.245 -11.395 ;
        RECT 393.555 -11.725 393.885 -11.395 ;
        RECT 392.195 -11.725 392.525 -11.395 ;
        RECT 390.835 -11.725 391.165 -11.395 ;
        RECT 389.475 -11.725 389.805 -11.395 ;
        RECT 388.115 -11.725 388.445 -11.395 ;
        RECT 386.755 -11.725 387.085 -11.395 ;
        RECT 385.395 -11.725 385.725 -11.395 ;
        RECT 384.035 -11.725 384.365 -11.395 ;
        RECT 382.675 -11.725 383.005 -11.395 ;
        RECT 381.315 -11.725 381.645 -11.395 ;
        RECT 379.955 -11.725 380.285 -11.395 ;
        RECT 378.595 -11.725 378.925 -11.395 ;
        RECT 377.235 -11.725 377.565 -11.395 ;
        RECT 375.875 -11.725 376.205 -11.395 ;
        RECT 374.515 -11.725 374.845 -11.395 ;
        RECT 373.155 -11.725 373.485 -11.395 ;
        RECT 371.795 -11.725 372.125 -11.395 ;
        RECT 370.435 -11.725 370.765 -11.395 ;
        RECT 369.075 -11.725 369.405 -11.395 ;
        RECT 367.715 -11.725 368.045 -11.395 ;
        RECT 366.355 -11.725 366.685 -11.395 ;
        RECT 364.995 -11.725 365.325 -11.395 ;
        RECT 363.635 -11.725 363.965 -11.395 ;
        RECT 362.275 -11.725 362.605 -11.395 ;
        RECT 360.915 -11.725 361.245 -11.395 ;
        RECT 359.555 -11.725 359.885 -11.395 ;
        RECT 358.195 -11.725 358.525 -11.395 ;
        RECT 356.835 -11.725 357.165 -11.395 ;
        RECT 355.475 -11.725 355.805 -11.395 ;
        RECT 354.115 -11.725 354.445 -11.395 ;
        RECT 352.755 -11.725 353.085 -11.395 ;
        RECT 351.395 -11.725 351.725 -11.395 ;
        RECT 350.035 -11.725 350.365 -11.395 ;
        RECT 348.675 -11.725 349.005 -11.395 ;
        RECT 347.315 -11.725 347.645 -11.395 ;
        RECT 345.955 -11.725 346.285 -11.395 ;
        RECT 344.595 -11.725 344.925 -11.395 ;
        RECT 343.235 -11.725 343.565 -11.395 ;
        RECT 341.875 -11.725 342.205 -11.395 ;
        RECT 340.515 -11.725 340.845 -11.395 ;
        RECT 339.155 -11.725 339.485 -11.395 ;
        RECT 337.795 -11.725 338.125 -11.395 ;
        RECT 336.435 -11.725 336.765 -11.395 ;
        RECT 335.075 -11.725 335.405 -11.395 ;
        RECT 333.715 -11.725 334.045 -11.395 ;
        RECT 332.355 -11.725 332.685 -11.395 ;
        RECT 330.995 -11.725 331.325 -11.395 ;
        RECT 329.635 -11.725 329.965 -11.395 ;
        RECT 328.275 -11.725 328.605 -11.395 ;
        RECT 326.915 -11.725 327.245 -11.395 ;
        RECT 325.555 -11.725 325.885 -11.395 ;
        RECT 324.195 -11.725 324.525 -11.395 ;
        RECT 322.835 -11.725 323.165 -11.395 ;
        RECT 321.475 -11.725 321.805 -11.395 ;
        RECT 320.115 -11.725 320.445 -11.395 ;
        RECT 318.755 -11.725 319.085 -11.395 ;
        RECT 317.395 -11.725 317.725 -11.395 ;
        RECT 316.035 -11.725 316.365 -11.395 ;
        RECT 314.675 -11.725 315.005 -11.395 ;
        RECT 313.315 -11.725 313.645 -11.395 ;
        RECT 311.955 -11.725 312.285 -11.395 ;
        RECT 310.595 -11.725 310.925 -11.395 ;
        RECT 309.235 -11.725 309.565 -11.395 ;
        RECT 307.875 -11.725 308.205 -11.395 ;
        RECT 306.515 -11.725 306.845 -11.395 ;
        RECT 305.155 -11.725 305.485 -11.395 ;
        RECT 303.795 -11.725 304.125 -11.395 ;
        RECT 302.435 -11.725 302.765 -11.395 ;
        RECT 301.075 -11.725 301.405 -11.395 ;
        RECT 299.715 -11.725 300.045 -11.395 ;
        RECT 298.355 -11.725 298.685 -11.395 ;
        RECT 296.995 -11.725 297.325 -11.395 ;
        RECT 295.635 -11.725 295.965 -11.395 ;
        RECT 294.275 -11.725 294.605 -11.395 ;
        RECT 292.915 -11.725 293.245 -11.395 ;
        RECT 291.555 -11.725 291.885 -11.395 ;
        RECT 290.195 -11.725 290.525 -11.395 ;
        RECT 288.835 -11.725 289.165 -11.395 ;
        RECT 287.475 -11.725 287.805 -11.395 ;
        RECT 286.115 -11.725 286.445 -11.395 ;
        RECT 284.755 -11.725 285.085 -11.395 ;
        RECT 283.395 -11.725 283.725 -11.395 ;
        RECT 282.035 -11.725 282.365 -11.395 ;
        RECT 280.675 -11.725 281.005 -11.395 ;
        RECT 279.315 -11.725 279.645 -11.395 ;
        RECT 277.955 -11.725 278.285 -11.395 ;
        RECT 276.595 -11.725 276.925 -11.395 ;
        RECT 275.235 -11.725 275.565 -11.395 ;
        RECT 273.875 -11.725 274.205 -11.395 ;
        RECT 272.515 -11.725 272.845 -11.395 ;
        RECT 271.155 -11.725 271.485 -11.395 ;
        RECT 269.795 -11.725 270.125 -11.395 ;
        RECT 268.435 -11.725 268.765 -11.395 ;
        RECT 267.075 -11.725 267.405 -11.395 ;
        RECT 265.715 -11.725 266.045 -11.395 ;
        RECT 264.355 -11.725 264.685 -11.395 ;
        RECT 262.995 -11.725 263.325 -11.395 ;
        RECT 261.635 -11.725 261.965 -11.395 ;
        RECT 260.275 -11.725 260.605 -11.395 ;
        RECT 258.915 -11.725 259.245 -11.395 ;
        RECT 257.555 -11.725 257.885 -11.395 ;
        RECT 256.195 -11.725 256.525 -11.395 ;
        RECT 254.835 -11.725 255.165 -11.395 ;
        RECT 253.475 -11.725 253.805 -11.395 ;
        RECT 252.115 -11.725 252.445 -11.395 ;
        RECT 250.755 -11.725 251.085 -11.395 ;
        RECT 249.395 -11.725 249.725 -11.395 ;
        RECT 248.035 -11.725 248.365 -11.395 ;
        RECT 246.675 -11.725 247.005 -11.395 ;
        RECT 245.315 -11.725 245.645 -11.395 ;
        RECT 243.955 -11.725 244.285 -11.395 ;
        RECT 242.595 -11.725 242.925 -11.395 ;
        RECT 241.235 -11.725 241.565 -11.395 ;
        RECT 239.875 -11.725 240.205 -11.395 ;
        RECT 238.515 -11.725 238.845 -11.395 ;
        RECT 237.155 -11.725 237.485 -11.395 ;
        RECT 235.795 -11.725 236.125 -11.395 ;
        RECT 234.435 -11.725 234.765 -11.395 ;
        RECT 233.075 -11.725 233.405 -11.395 ;
        RECT 231.715 -11.725 232.045 -11.395 ;
        RECT 230.355 -11.725 230.685 -11.395 ;
        RECT 228.995 -11.725 229.325 -11.395 ;
        RECT 227.635 -11.725 227.965 -11.395 ;
        RECT 226.275 -11.725 226.605 -11.395 ;
        RECT 224.915 -11.725 225.245 -11.395 ;
        RECT 223.555 -11.725 223.885 -11.395 ;
        RECT 222.195 -11.725 222.525 -11.395 ;
        RECT 220.835 -11.725 221.165 -11.395 ;
        RECT 219.475 -11.725 219.805 -11.395 ;
        RECT 218.115 -11.725 218.445 -11.395 ;
        RECT 216.755 -11.725 217.085 -11.395 ;
        RECT 215.395 -11.725 215.725 -11.395 ;
        RECT 214.035 -11.725 214.365 -11.395 ;
        RECT 212.675 -11.725 213.005 -11.395 ;
        RECT 211.315 -11.725 211.645 -11.395 ;
        RECT 209.955 -11.725 210.285 -11.395 ;
        RECT 208.595 -11.725 208.925 -11.395 ;
        RECT 207.235 -11.725 207.565 -11.395 ;
        RECT 205.875 -11.725 206.205 -11.395 ;
        RECT 204.515 -11.725 204.845 -11.395 ;
        RECT 203.155 -11.725 203.485 -11.395 ;
        RECT 201.795 -11.725 202.125 -11.395 ;
        RECT 200.435 -11.725 200.765 -11.395 ;
        RECT 199.075 -11.725 199.405 -11.395 ;
        RECT 197.715 -11.725 198.045 -11.395 ;
        RECT 196.355 -11.725 196.685 -11.395 ;
        RECT 194.995 -11.725 195.325 -11.395 ;
        RECT 193.635 -11.725 193.965 -11.395 ;
        RECT 192.275 -11.725 192.605 -11.395 ;
        RECT 190.915 -11.725 191.245 -11.395 ;
        RECT 189.555 -11.725 189.885 -11.395 ;
        RECT 188.195 -11.725 188.525 -11.395 ;
        RECT 186.835 -11.725 187.165 -11.395 ;
        RECT 185.475 -11.725 185.805 -11.395 ;
        RECT 184.115 -11.725 184.445 -11.395 ;
        RECT 182.755 -11.725 183.085 -11.395 ;
        RECT 181.395 -11.725 181.725 -11.395 ;
        RECT 180.035 -11.725 180.365 -11.395 ;
        RECT 178.675 -11.725 179.005 -11.395 ;
        RECT 177.315 -11.725 177.645 -11.395 ;
        RECT 175.955 -11.725 176.285 -11.395 ;
        RECT 174.595 -11.725 174.925 -11.395 ;
        RECT 173.235 -11.725 173.565 -11.395 ;
        RECT 171.875 -11.725 172.205 -11.395 ;
        RECT 170.515 -11.725 170.845 -11.395 ;
        RECT 169.155 -11.725 169.485 -11.395 ;
        RECT 167.795 -11.725 168.125 -11.395 ;
        RECT 166.435 -11.725 166.765 -11.395 ;
        RECT 165.075 -11.725 165.405 -11.395 ;
        RECT 163.715 -11.725 164.045 -11.395 ;
        RECT 162.355 -11.725 162.685 -11.395 ;
        RECT 160.995 -11.725 161.325 -11.395 ;
        RECT 159.635 -11.725 159.965 -11.395 ;
        RECT 158.275 -11.725 158.605 -11.395 ;
        RECT 156.915 -11.725 157.245 -11.395 ;
        RECT 155.555 -11.725 155.885 -11.395 ;
        RECT 154.195 -11.725 154.525 -11.395 ;
        RECT 152.835 -11.725 153.165 -11.395 ;
        RECT 151.475 -11.725 151.805 -11.395 ;
        RECT 150.115 -11.725 150.445 -11.395 ;
        RECT 148.755 -11.725 149.085 -11.395 ;
        RECT 147.395 -11.725 147.725 -11.395 ;
        RECT 146.035 -11.725 146.365 -11.395 ;
        RECT 144.675 -11.725 145.005 -11.395 ;
        RECT 143.315 -11.725 143.645 -11.395 ;
        RECT 141.955 -11.725 142.285 -11.395 ;
        RECT 140.595 -11.725 140.925 -11.395 ;
        RECT 139.235 -11.725 139.565 -11.395 ;
        RECT 137.875 -11.725 138.205 -11.395 ;
        RECT 136.515 -11.725 136.845 -11.395 ;
        RECT 135.155 -11.725 135.485 -11.395 ;
        RECT 133.795 -11.725 134.125 -11.395 ;
        RECT 132.435 -11.725 132.765 -11.395 ;
        RECT 131.075 -11.725 131.405 -11.395 ;
        RECT 129.715 -11.725 130.045 -11.395 ;
        RECT 734.915 -11.725 735.245 -11.395 ;
        RECT 733.555 -11.725 733.885 -11.395 ;
        RECT 732.195 -11.725 732.525 -11.395 ;
        RECT 730.835 -11.725 731.165 -11.395 ;
        RECT 729.475 -11.725 729.805 -11.395 ;
        RECT 728.115 -11.725 728.445 -11.395 ;
        RECT 726.755 -11.725 727.085 -11.395 ;
        RECT 725.395 -11.725 725.725 -11.395 ;
        RECT 724.035 -11.725 724.365 -11.395 ;
        RECT 722.675 -11.725 723.005 -11.395 ;
        RECT 721.315 -11.725 721.645 -11.395 ;
        RECT 719.955 -11.725 720.285 -11.395 ;
        RECT 718.595 -11.725 718.925 -11.395 ;
        RECT 717.235 -11.725 717.565 -11.395 ;
        RECT 715.875 -11.725 716.205 -11.395 ;
        RECT 714.515 -11.725 714.845 -11.395 ;
        RECT 713.155 -11.725 713.485 -11.395 ;
        RECT 711.795 -11.725 712.125 -11.395 ;
        RECT 710.435 -11.725 710.765 -11.395 ;
        RECT 709.075 -11.725 709.405 -11.395 ;
        RECT 707.715 -11.725 708.045 -11.395 ;
        RECT 706.355 -11.725 706.685 -11.395 ;
        RECT 704.995 -11.725 705.325 -11.395 ;
        RECT 703.635 -11.725 703.965 -11.395 ;
        RECT 702.275 -11.725 702.605 -11.395 ;
        RECT 700.915 -11.725 701.245 -11.395 ;
        RECT 699.555 -11.725 699.885 -11.395 ;
        RECT 698.195 -11.725 698.525 -11.395 ;
        RECT 696.835 -11.725 697.165 -11.395 ;
        RECT 695.475 -11.725 695.805 -11.395 ;
        RECT 694.115 -11.725 694.445 -11.395 ;
        RECT 692.755 -11.725 693.085 -11.395 ;
        RECT 691.395 -11.725 691.725 -11.395 ;
        RECT 690.035 -11.725 690.365 -11.395 ;
        RECT 688.675 -11.725 689.005 -11.395 ;
        RECT 687.315 -11.725 687.645 -11.395 ;
        RECT 685.955 -11.725 686.285 -11.395 ;
        RECT 684.595 -11.725 684.925 -11.395 ;
        RECT 683.235 -11.725 683.565 -11.395 ;
        RECT 681.875 -11.725 682.205 -11.395 ;
        RECT 680.515 -11.725 680.845 -11.395 ;
        RECT 679.155 -11.725 679.485 -11.395 ;
        RECT 678.125 -11.72 954.88 -11.4 ;
        RECT 953.875 -11.725 954.205 -11.395 ;
        RECT 952.515 -11.725 952.845 -11.395 ;
        RECT 951.155 -11.725 951.485 -11.395 ;
        RECT 949.795 -11.725 950.125 -11.395 ;
        RECT 948.435 -11.725 948.765 -11.395 ;
        RECT 947.075 -11.725 947.405 -11.395 ;
        RECT 945.715 -11.725 946.045 -11.395 ;
        RECT 944.355 -11.725 944.685 -11.395 ;
        RECT 942.995 -11.725 943.325 -11.395 ;
        RECT 941.635 -11.725 941.965 -11.395 ;
        RECT 940.275 -11.725 940.605 -11.395 ;
        RECT 938.915 -11.725 939.245 -11.395 ;
        RECT 937.555 -11.725 937.885 -11.395 ;
        RECT 936.195 -11.725 936.525 -11.395 ;
        RECT 934.835 -11.725 935.165 -11.395 ;
        RECT 933.475 -11.725 933.805 -11.395 ;
        RECT 932.115 -11.725 932.445 -11.395 ;
        RECT 930.755 -11.725 931.085 -11.395 ;
        RECT 929.395 -11.725 929.725 -11.395 ;
        RECT 928.035 -11.725 928.365 -11.395 ;
        RECT 926.675 -11.725 927.005 -11.395 ;
        RECT 925.315 -11.725 925.645 -11.395 ;
        RECT 923.955 -11.725 924.285 -11.395 ;
        RECT 922.595 -11.725 922.925 -11.395 ;
        RECT 921.235 -11.725 921.565 -11.395 ;
        RECT 919.875 -11.725 920.205 -11.395 ;
        RECT 918.515 -11.725 918.845 -11.395 ;
        RECT 917.155 -11.725 917.485 -11.395 ;
        RECT 915.795 -11.725 916.125 -11.395 ;
        RECT 914.435 -11.725 914.765 -11.395 ;
        RECT 913.075 -11.725 913.405 -11.395 ;
        RECT 911.715 -11.725 912.045 -11.395 ;
        RECT 910.355 -11.725 910.685 -11.395 ;
        RECT 908.995 -11.725 909.325 -11.395 ;
        RECT 907.635 -11.725 907.965 -11.395 ;
        RECT 906.275 -11.725 906.605 -11.395 ;
        RECT 904.915 -11.725 905.245 -11.395 ;
        RECT 903.555 -11.725 903.885 -11.395 ;
        RECT 902.195 -11.725 902.525 -11.395 ;
        RECT 900.835 -11.725 901.165 -11.395 ;
        RECT 899.475 -11.725 899.805 -11.395 ;
        RECT 898.115 -11.725 898.445 -11.395 ;
        RECT 896.755 -11.725 897.085 -11.395 ;
        RECT 895.395 -11.725 895.725 -11.395 ;
        RECT 894.035 -11.725 894.365 -11.395 ;
        RECT 892.675 -11.725 893.005 -11.395 ;
        RECT 891.315 -11.725 891.645 -11.395 ;
        RECT 889.955 -11.725 890.285 -11.395 ;
        RECT 888.595 -11.725 888.925 -11.395 ;
        RECT 887.235 -11.725 887.565 -11.395 ;
        RECT 885.875 -11.725 886.205 -11.395 ;
        RECT 884.515 -11.725 884.845 -11.395 ;
        RECT 883.155 -11.725 883.485 -11.395 ;
        RECT 881.795 -11.725 882.125 -11.395 ;
        RECT 880.435 -11.725 880.765 -11.395 ;
        RECT 879.075 -11.725 879.405 -11.395 ;
        RECT 877.715 -11.725 878.045 -11.395 ;
        RECT 876.355 -11.725 876.685 -11.395 ;
        RECT 874.995 -11.725 875.325 -11.395 ;
        RECT 873.635 -11.725 873.965 -11.395 ;
        RECT 872.275 -11.725 872.605 -11.395 ;
        RECT 870.915 -11.725 871.245 -11.395 ;
        RECT 869.555 -11.725 869.885 -11.395 ;
        RECT 868.195 -11.725 868.525 -11.395 ;
        RECT 866.835 -11.725 867.165 -11.395 ;
        RECT 865.475 -11.725 865.805 -11.395 ;
        RECT 864.115 -11.725 864.445 -11.395 ;
        RECT 862.755 -11.725 863.085 -11.395 ;
        RECT 861.395 -11.725 861.725 -11.395 ;
        RECT 860.035 -11.725 860.365 -11.395 ;
        RECT 858.675 -11.725 859.005 -11.395 ;
        RECT 857.315 -11.725 857.645 -11.395 ;
        RECT 855.955 -11.725 856.285 -11.395 ;
        RECT 854.595 -11.725 854.925 -11.395 ;
        RECT 853.235 -11.725 853.565 -11.395 ;
        RECT 851.875 -11.725 852.205 -11.395 ;
        RECT 850.515 -11.725 850.845 -11.395 ;
        RECT 849.155 -11.725 849.485 -11.395 ;
        RECT 847.795 -11.725 848.125 -11.395 ;
        RECT 846.435 -11.725 846.765 -11.395 ;
        RECT 845.075 -11.725 845.405 -11.395 ;
        RECT 843.715 -11.725 844.045 -11.395 ;
        RECT 842.355 -11.725 842.685 -11.395 ;
        RECT 840.995 -11.725 841.325 -11.395 ;
        RECT 839.635 -11.725 839.965 -11.395 ;
        RECT 838.275 -11.725 838.605 -11.395 ;
        RECT 836.915 -11.725 837.245 -11.395 ;
        RECT 835.555 -11.725 835.885 -11.395 ;
        RECT 834.195 -11.725 834.525 -11.395 ;
        RECT 832.835 -11.725 833.165 -11.395 ;
        RECT 831.475 -11.725 831.805 -11.395 ;
        RECT 830.115 -11.725 830.445 -11.395 ;
        RECT 828.755 -11.725 829.085 -11.395 ;
        RECT 827.395 -11.725 827.725 -11.395 ;
        RECT 826.035 -11.725 826.365 -11.395 ;
        RECT 824.675 -11.725 825.005 -11.395 ;
        RECT 823.315 -11.725 823.645 -11.395 ;
        RECT 821.955 -11.725 822.285 -11.395 ;
        RECT 820.595 -11.725 820.925 -11.395 ;
        RECT 819.235 -11.725 819.565 -11.395 ;
        RECT 817.875 -11.725 818.205 -11.395 ;
        RECT 816.515 -11.725 816.845 -11.395 ;
        RECT 815.155 -11.725 815.485 -11.395 ;
        RECT 813.795 -11.725 814.125 -11.395 ;
        RECT 812.435 -11.725 812.765 -11.395 ;
        RECT 811.075 -11.725 811.405 -11.395 ;
        RECT 809.715 -11.725 810.045 -11.395 ;
        RECT 808.355 -11.725 808.685 -11.395 ;
        RECT 806.995 -11.725 807.325 -11.395 ;
        RECT 805.635 -11.725 805.965 -11.395 ;
        RECT 804.275 -11.725 804.605 -11.395 ;
        RECT 802.915 -11.725 803.245 -11.395 ;
        RECT 801.555 -11.725 801.885 -11.395 ;
        RECT 800.195 -11.725 800.525 -11.395 ;
        RECT 798.835 -11.725 799.165 -11.395 ;
        RECT 797.475 -11.725 797.805 -11.395 ;
        RECT 796.115 -11.725 796.445 -11.395 ;
        RECT 794.755 -11.725 795.085 -11.395 ;
        RECT 793.395 -11.725 793.725 -11.395 ;
        RECT 792.035 -11.725 792.365 -11.395 ;
        RECT 790.675 -11.725 791.005 -11.395 ;
        RECT 789.315 -11.725 789.645 -11.395 ;
        RECT 787.955 -11.725 788.285 -11.395 ;
        RECT 786.595 -11.725 786.925 -11.395 ;
        RECT 785.235 -11.725 785.565 -11.395 ;
        RECT 783.875 -11.725 784.205 -11.395 ;
        RECT 782.515 -11.725 782.845 -11.395 ;
        RECT 781.155 -11.725 781.485 -11.395 ;
        RECT 779.795 -11.725 780.125 -11.395 ;
        RECT 778.435 -11.725 778.765 -11.395 ;
        RECT 777.075 -11.725 777.405 -11.395 ;
        RECT 775.715 -11.725 776.045 -11.395 ;
        RECT 774.355 -11.725 774.685 -11.395 ;
        RECT 772.995 -11.725 773.325 -11.395 ;
        RECT 771.635 -11.725 771.965 -11.395 ;
        RECT 770.275 -11.725 770.605 -11.395 ;
        RECT 768.915 -11.725 769.245 -11.395 ;
        RECT 767.555 -11.725 767.885 -11.395 ;
        RECT 766.195 -11.725 766.525 -11.395 ;
        RECT 764.835 -11.725 765.165 -11.395 ;
        RECT 763.475 -11.725 763.805 -11.395 ;
        RECT 762.115 -11.725 762.445 -11.395 ;
        RECT 760.755 -11.725 761.085 -11.395 ;
        RECT 759.395 -11.725 759.725 -11.395 ;
        RECT 758.035 -11.725 758.365 -11.395 ;
        RECT 756.675 -11.725 757.005 -11.395 ;
        RECT 755.315 -11.725 755.645 -11.395 ;
        RECT 753.955 -11.725 754.285 -11.395 ;
        RECT 752.595 -11.725 752.925 -11.395 ;
        RECT 751.235 -11.725 751.565 -11.395 ;
        RECT 749.875 -11.725 750.205 -11.395 ;
        RECT 748.515 -11.725 748.845 -11.395 ;
        RECT 747.155 -11.725 747.485 -11.395 ;
        RECT 745.795 -11.725 746.125 -11.395 ;
        RECT 744.435 -11.725 744.765 -11.395 ;
        RECT 743.075 -11.725 743.405 -11.395 ;
        RECT 741.715 -11.725 742.045 -11.395 ;
        RECT 740.355 -11.725 740.685 -11.395 ;
        RECT 738.995 -11.725 739.325 -11.395 ;
        RECT 737.635 -11.725 737.965 -11.395 ;
        RECT 736.275 -11.725 736.605 -11.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 -7.645 678.125 -7.315 ;
        RECT -1.52 -7.64 678.125 -7.32 ;
        RECT 676.435 -7.645 676.765 -7.315 ;
        RECT 675.075 -7.645 675.405 -7.315 ;
        RECT 673.715 -7.645 674.045 -7.315 ;
        RECT 672.355 -7.645 672.685 -7.315 ;
        RECT 670.995 -7.645 671.325 -7.315 ;
        RECT 669.635 -7.645 669.965 -7.315 ;
        RECT 668.275 -7.645 668.605 -7.315 ;
        RECT 666.915 -7.645 667.245 -7.315 ;
        RECT 665.555 -7.645 665.885 -7.315 ;
        RECT 664.195 -7.645 664.525 -7.315 ;
        RECT 662.835 -7.645 663.165 -7.315 ;
        RECT 661.475 -7.645 661.805 -7.315 ;
        RECT 660.115 -7.645 660.445 -7.315 ;
        RECT 658.755 -7.645 659.085 -7.315 ;
        RECT 657.395 -7.645 657.725 -7.315 ;
        RECT 656.035 -7.645 656.365 -7.315 ;
        RECT 654.675 -7.645 655.005 -7.315 ;
        RECT 653.315 -7.645 653.645 -7.315 ;
        RECT 651.955 -7.645 652.285 -7.315 ;
        RECT 650.595 -7.645 650.925 -7.315 ;
        RECT 649.235 -7.645 649.565 -7.315 ;
        RECT 647.875 -7.645 648.205 -7.315 ;
        RECT 646.515 -7.645 646.845 -7.315 ;
        RECT 645.155 -7.645 645.485 -7.315 ;
        RECT 643.795 -7.645 644.125 -7.315 ;
        RECT 642.435 -7.645 642.765 -7.315 ;
        RECT 641.075 -7.645 641.405 -7.315 ;
        RECT 639.715 -7.645 640.045 -7.315 ;
        RECT 638.355 -7.645 638.685 -7.315 ;
        RECT 636.995 -7.645 637.325 -7.315 ;
        RECT 635.635 -7.645 635.965 -7.315 ;
        RECT 634.275 -7.645 634.605 -7.315 ;
        RECT 632.915 -7.645 633.245 -7.315 ;
        RECT 631.555 -7.645 631.885 -7.315 ;
        RECT 630.195 -7.645 630.525 -7.315 ;
        RECT 628.835 -7.645 629.165 -7.315 ;
        RECT 627.475 -7.645 627.805 -7.315 ;
        RECT 626.115 -7.645 626.445 -7.315 ;
        RECT 624.755 -7.645 625.085 -7.315 ;
        RECT 623.395 -7.645 623.725 -7.315 ;
        RECT 622.035 -7.645 622.365 -7.315 ;
        RECT 620.675 -7.645 621.005 -7.315 ;
        RECT 619.315 -7.645 619.645 -7.315 ;
        RECT 617.955 -7.645 618.285 -7.315 ;
        RECT 616.595 -7.645 616.925 -7.315 ;
        RECT 615.235 -7.645 615.565 -7.315 ;
        RECT 613.875 -7.645 614.205 -7.315 ;
        RECT 612.515 -7.645 612.845 -7.315 ;
        RECT 611.155 -7.645 611.485 -7.315 ;
        RECT 609.795 -7.645 610.125 -7.315 ;
        RECT 608.435 -7.645 608.765 -7.315 ;
        RECT 607.075 -7.645 607.405 -7.315 ;
        RECT 605.715 -7.645 606.045 -7.315 ;
        RECT 604.355 -7.645 604.685 -7.315 ;
        RECT 602.995 -7.645 603.325 -7.315 ;
        RECT 601.635 -7.645 601.965 -7.315 ;
        RECT 600.275 -7.645 600.605 -7.315 ;
        RECT 598.915 -7.645 599.245 -7.315 ;
        RECT 597.555 -7.645 597.885 -7.315 ;
        RECT 596.195 -7.645 596.525 -7.315 ;
        RECT 594.835 -7.645 595.165 -7.315 ;
        RECT 593.475 -7.645 593.805 -7.315 ;
        RECT 592.115 -7.645 592.445 -7.315 ;
        RECT 590.755 -7.645 591.085 -7.315 ;
        RECT 589.395 -7.645 589.725 -7.315 ;
        RECT 588.035 -7.645 588.365 -7.315 ;
        RECT 586.675 -7.645 587.005 -7.315 ;
        RECT 585.315 -7.645 585.645 -7.315 ;
        RECT 583.955 -7.645 584.285 -7.315 ;
        RECT 582.595 -7.645 582.925 -7.315 ;
        RECT 581.235 -7.645 581.565 -7.315 ;
        RECT 579.875 -7.645 580.205 -7.315 ;
        RECT 578.515 -7.645 578.845 -7.315 ;
        RECT 577.155 -7.645 577.485 -7.315 ;
        RECT 575.795 -7.645 576.125 -7.315 ;
        RECT 574.435 -7.645 574.765 -7.315 ;
        RECT 573.075 -7.645 573.405 -7.315 ;
        RECT 571.715 -7.645 572.045 -7.315 ;
        RECT 570.355 -7.645 570.685 -7.315 ;
        RECT 568.995 -7.645 569.325 -7.315 ;
        RECT 567.635 -7.645 567.965 -7.315 ;
        RECT 566.275 -7.645 566.605 -7.315 ;
        RECT 564.915 -7.645 565.245 -7.315 ;
        RECT 563.555 -7.645 563.885 -7.315 ;
        RECT 562.195 -7.645 562.525 -7.315 ;
        RECT 560.835 -7.645 561.165 -7.315 ;
        RECT 559.475 -7.645 559.805 -7.315 ;
        RECT 558.115 -7.645 558.445 -7.315 ;
        RECT 556.755 -7.645 557.085 -7.315 ;
        RECT 555.395 -7.645 555.725 -7.315 ;
        RECT 554.035 -7.645 554.365 -7.315 ;
        RECT 552.675 -7.645 553.005 -7.315 ;
        RECT 551.315 -7.645 551.645 -7.315 ;
        RECT 549.955 -7.645 550.285 -7.315 ;
        RECT 548.595 -7.645 548.925 -7.315 ;
        RECT 547.235 -7.645 547.565 -7.315 ;
        RECT 545.875 -7.645 546.205 -7.315 ;
        RECT 544.515 -7.645 544.845 -7.315 ;
        RECT 543.155 -7.645 543.485 -7.315 ;
        RECT 541.795 -7.645 542.125 -7.315 ;
        RECT 540.435 -7.645 540.765 -7.315 ;
        RECT 539.075 -7.645 539.405 -7.315 ;
        RECT 537.715 -7.645 538.045 -7.315 ;
        RECT 536.355 -7.645 536.685 -7.315 ;
        RECT 534.995 -7.645 535.325 -7.315 ;
        RECT 533.635 -7.645 533.965 -7.315 ;
        RECT 532.275 -7.645 532.605 -7.315 ;
        RECT 530.915 -7.645 531.245 -7.315 ;
        RECT 529.555 -7.645 529.885 -7.315 ;
        RECT 528.195 -7.645 528.525 -7.315 ;
        RECT 526.835 -7.645 527.165 -7.315 ;
        RECT 525.475 -7.645 525.805 -7.315 ;
        RECT 524.115 -7.645 524.445 -7.315 ;
        RECT 522.755 -7.645 523.085 -7.315 ;
        RECT 521.395 -7.645 521.725 -7.315 ;
        RECT 520.035 -7.645 520.365 -7.315 ;
        RECT 518.675 -7.645 519.005 -7.315 ;
        RECT 517.315 -7.645 517.645 -7.315 ;
        RECT 515.955 -7.645 516.285 -7.315 ;
        RECT 514.595 -7.645 514.925 -7.315 ;
        RECT 513.235 -7.645 513.565 -7.315 ;
        RECT 511.875 -7.645 512.205 -7.315 ;
        RECT 510.515 -7.645 510.845 -7.315 ;
        RECT 509.155 -7.645 509.485 -7.315 ;
        RECT 507.795 -7.645 508.125 -7.315 ;
        RECT 506.435 -7.645 506.765 -7.315 ;
        RECT 505.075 -7.645 505.405 -7.315 ;
        RECT 503.715 -7.645 504.045 -7.315 ;
        RECT 502.355 -7.645 502.685 -7.315 ;
        RECT 500.995 -7.645 501.325 -7.315 ;
        RECT 499.635 -7.645 499.965 -7.315 ;
        RECT 498.275 -7.645 498.605 -7.315 ;
        RECT 496.915 -7.645 497.245 -7.315 ;
        RECT 495.555 -7.645 495.885 -7.315 ;
        RECT 494.195 -7.645 494.525 -7.315 ;
        RECT 492.835 -7.645 493.165 -7.315 ;
        RECT 491.475 -7.645 491.805 -7.315 ;
        RECT 490.115 -7.645 490.445 -7.315 ;
        RECT 488.755 -7.645 489.085 -7.315 ;
        RECT 487.395 -7.645 487.725 -7.315 ;
        RECT 486.035 -7.645 486.365 -7.315 ;
        RECT 484.675 -7.645 485.005 -7.315 ;
        RECT 483.315 -7.645 483.645 -7.315 ;
        RECT 481.955 -7.645 482.285 -7.315 ;
        RECT 480.595 -7.645 480.925 -7.315 ;
        RECT 479.235 -7.645 479.565 -7.315 ;
        RECT 477.875 -7.645 478.205 -7.315 ;
        RECT 476.515 -7.645 476.845 -7.315 ;
        RECT 475.155 -7.645 475.485 -7.315 ;
        RECT 473.795 -7.645 474.125 -7.315 ;
        RECT 472.435 -7.645 472.765 -7.315 ;
        RECT 471.075 -7.645 471.405 -7.315 ;
        RECT 469.715 -7.645 470.045 -7.315 ;
        RECT 468.355 -7.645 468.685 -7.315 ;
        RECT 466.995 -7.645 467.325 -7.315 ;
        RECT 465.635 -7.645 465.965 -7.315 ;
        RECT 464.275 -7.645 464.605 -7.315 ;
        RECT 462.915 -7.645 463.245 -7.315 ;
        RECT 461.555 -7.645 461.885 -7.315 ;
        RECT 460.195 -7.645 460.525 -7.315 ;
        RECT 458.835 -7.645 459.165 -7.315 ;
        RECT 457.475 -7.645 457.805 -7.315 ;
        RECT 456.115 -7.645 456.445 -7.315 ;
        RECT 454.755 -7.645 455.085 -7.315 ;
        RECT 453.395 -7.645 453.725 -7.315 ;
        RECT 452.035 -7.645 452.365 -7.315 ;
        RECT 450.675 -7.645 451.005 -7.315 ;
        RECT 449.315 -7.645 449.645 -7.315 ;
        RECT 447.955 -7.645 448.285 -7.315 ;
        RECT 446.595 -7.645 446.925 -7.315 ;
        RECT 445.235 -7.645 445.565 -7.315 ;
        RECT 443.875 -7.645 444.205 -7.315 ;
        RECT 442.515 -7.645 442.845 -7.315 ;
        RECT 441.155 -7.645 441.485 -7.315 ;
        RECT 439.795 -7.645 440.125 -7.315 ;
        RECT 438.435 -7.645 438.765 -7.315 ;
        RECT 437.075 -7.645 437.405 -7.315 ;
        RECT 435.715 -7.645 436.045 -7.315 ;
        RECT 434.355 -7.645 434.685 -7.315 ;
        RECT 432.995 -7.645 433.325 -7.315 ;
        RECT 431.635 -7.645 431.965 -7.315 ;
        RECT 430.275 -7.645 430.605 -7.315 ;
        RECT 428.915 -7.645 429.245 -7.315 ;
        RECT 427.555 -7.645 427.885 -7.315 ;
        RECT 426.195 -7.645 426.525 -7.315 ;
        RECT 424.835 -7.645 425.165 -7.315 ;
        RECT 423.475 -7.645 423.805 -7.315 ;
        RECT 422.115 -7.645 422.445 -7.315 ;
        RECT 420.755 -7.645 421.085 -7.315 ;
        RECT 419.395 -7.645 419.725 -7.315 ;
        RECT 418.035 -7.645 418.365 -7.315 ;
        RECT 416.675 -7.645 417.005 -7.315 ;
        RECT 415.315 -7.645 415.645 -7.315 ;
        RECT 413.955 -7.645 414.285 -7.315 ;
        RECT 412.595 -7.645 412.925 -7.315 ;
        RECT 411.235 -7.645 411.565 -7.315 ;
        RECT 409.875 -7.645 410.205 -7.315 ;
        RECT 408.515 -7.645 408.845 -7.315 ;
        RECT 407.155 -7.645 407.485 -7.315 ;
        RECT 405.795 -7.645 406.125 -7.315 ;
        RECT 404.435 -7.645 404.765 -7.315 ;
        RECT 403.075 -7.645 403.405 -7.315 ;
        RECT 401.715 -7.645 402.045 -7.315 ;
        RECT 400.355 -7.645 400.685 -7.315 ;
        RECT 398.995 -7.645 399.325 -7.315 ;
        RECT 397.635 -7.645 397.965 -7.315 ;
        RECT 396.275 -7.645 396.605 -7.315 ;
        RECT 394.915 -7.645 395.245 -7.315 ;
        RECT 393.555 -7.645 393.885 -7.315 ;
        RECT 392.195 -7.645 392.525 -7.315 ;
        RECT 390.835 -7.645 391.165 -7.315 ;
        RECT 389.475 -7.645 389.805 -7.315 ;
        RECT 388.115 -7.645 388.445 -7.315 ;
        RECT 386.755 -7.645 387.085 -7.315 ;
        RECT 385.395 -7.645 385.725 -7.315 ;
        RECT 384.035 -7.645 384.365 -7.315 ;
        RECT 382.675 -7.645 383.005 -7.315 ;
        RECT 381.315 -7.645 381.645 -7.315 ;
        RECT 379.955 -7.645 380.285 -7.315 ;
        RECT 378.595 -7.645 378.925 -7.315 ;
        RECT 377.235 -7.645 377.565 -7.315 ;
        RECT 375.875 -7.645 376.205 -7.315 ;
        RECT 374.515 -7.645 374.845 -7.315 ;
        RECT 373.155 -7.645 373.485 -7.315 ;
        RECT 371.795 -7.645 372.125 -7.315 ;
        RECT 370.435 -7.645 370.765 -7.315 ;
        RECT 369.075 -7.645 369.405 -7.315 ;
        RECT 367.715 -7.645 368.045 -7.315 ;
        RECT 366.355 -7.645 366.685 -7.315 ;
        RECT 364.995 -7.645 365.325 -7.315 ;
        RECT 363.635 -7.645 363.965 -7.315 ;
        RECT 362.275 -7.645 362.605 -7.315 ;
        RECT 360.915 -7.645 361.245 -7.315 ;
        RECT 359.555 -7.645 359.885 -7.315 ;
        RECT 358.195 -7.645 358.525 -7.315 ;
        RECT 356.835 -7.645 357.165 -7.315 ;
        RECT 355.475 -7.645 355.805 -7.315 ;
        RECT 354.115 -7.645 354.445 -7.315 ;
        RECT 352.755 -7.645 353.085 -7.315 ;
        RECT 351.395 -7.645 351.725 -7.315 ;
        RECT 350.035 -7.645 350.365 -7.315 ;
        RECT 348.675 -7.645 349.005 -7.315 ;
        RECT 347.315 -7.645 347.645 -7.315 ;
        RECT 345.955 -7.645 346.285 -7.315 ;
        RECT 344.595 -7.645 344.925 -7.315 ;
        RECT 343.235 -7.645 343.565 -7.315 ;
        RECT 341.875 -7.645 342.205 -7.315 ;
        RECT 340.515 -7.645 340.845 -7.315 ;
        RECT 339.155 -7.645 339.485 -7.315 ;
        RECT 337.795 -7.645 338.125 -7.315 ;
        RECT 336.435 -7.645 336.765 -7.315 ;
        RECT 335.075 -7.645 335.405 -7.315 ;
        RECT 333.715 -7.645 334.045 -7.315 ;
        RECT 332.355 -7.645 332.685 -7.315 ;
        RECT 330.995 -7.645 331.325 -7.315 ;
        RECT 329.635 -7.645 329.965 -7.315 ;
        RECT 328.275 -7.645 328.605 -7.315 ;
        RECT 326.915 -7.645 327.245 -7.315 ;
        RECT 325.555 -7.645 325.885 -7.315 ;
        RECT 324.195 -7.645 324.525 -7.315 ;
        RECT 322.835 -7.645 323.165 -7.315 ;
        RECT 321.475 -7.645 321.805 -7.315 ;
        RECT 320.115 -7.645 320.445 -7.315 ;
        RECT 318.755 -7.645 319.085 -7.315 ;
        RECT 317.395 -7.645 317.725 -7.315 ;
        RECT 316.035 -7.645 316.365 -7.315 ;
        RECT 314.675 -7.645 315.005 -7.315 ;
        RECT 313.315 -7.645 313.645 -7.315 ;
        RECT 311.955 -7.645 312.285 -7.315 ;
        RECT 310.595 -7.645 310.925 -7.315 ;
        RECT 309.235 -7.645 309.565 -7.315 ;
        RECT 307.875 -7.645 308.205 -7.315 ;
        RECT 306.515 -7.645 306.845 -7.315 ;
        RECT 305.155 -7.645 305.485 -7.315 ;
        RECT 303.795 -7.645 304.125 -7.315 ;
        RECT 302.435 -7.645 302.765 -7.315 ;
        RECT 301.075 -7.645 301.405 -7.315 ;
        RECT 299.715 -7.645 300.045 -7.315 ;
        RECT 298.355 -7.645 298.685 -7.315 ;
        RECT 296.995 -7.645 297.325 -7.315 ;
        RECT 295.635 -7.645 295.965 -7.315 ;
        RECT 294.275 -7.645 294.605 -7.315 ;
        RECT 292.915 -7.645 293.245 -7.315 ;
        RECT 291.555 -7.645 291.885 -7.315 ;
        RECT 290.195 -7.645 290.525 -7.315 ;
        RECT 288.835 -7.645 289.165 -7.315 ;
        RECT 287.475 -7.645 287.805 -7.315 ;
        RECT 286.115 -7.645 286.445 -7.315 ;
        RECT 284.755 -7.645 285.085 -7.315 ;
        RECT 283.395 -7.645 283.725 -7.315 ;
        RECT 282.035 -7.645 282.365 -7.315 ;
        RECT 280.675 -7.645 281.005 -7.315 ;
        RECT 279.315 -7.645 279.645 -7.315 ;
        RECT 277.955 -7.645 278.285 -7.315 ;
        RECT 276.595 -7.645 276.925 -7.315 ;
        RECT 275.235 -7.645 275.565 -7.315 ;
        RECT 273.875 -7.645 274.205 -7.315 ;
        RECT 272.515 -7.645 272.845 -7.315 ;
        RECT 271.155 -7.645 271.485 -7.315 ;
        RECT 269.795 -7.645 270.125 -7.315 ;
        RECT 268.435 -7.645 268.765 -7.315 ;
        RECT 267.075 -7.645 267.405 -7.315 ;
        RECT 265.715 -7.645 266.045 -7.315 ;
        RECT 264.355 -7.645 264.685 -7.315 ;
        RECT 262.995 -7.645 263.325 -7.315 ;
        RECT 261.635 -7.645 261.965 -7.315 ;
        RECT 260.275 -7.645 260.605 -7.315 ;
        RECT 258.915 -7.645 259.245 -7.315 ;
        RECT 257.555 -7.645 257.885 -7.315 ;
        RECT 256.195 -7.645 256.525 -7.315 ;
        RECT 254.835 -7.645 255.165 -7.315 ;
        RECT 253.475 -7.645 253.805 -7.315 ;
        RECT 252.115 -7.645 252.445 -7.315 ;
        RECT 250.755 -7.645 251.085 -7.315 ;
        RECT 249.395 -7.645 249.725 -7.315 ;
        RECT 248.035 -7.645 248.365 -7.315 ;
        RECT 246.675 -7.645 247.005 -7.315 ;
        RECT 245.315 -7.645 245.645 -7.315 ;
        RECT 243.955 -7.645 244.285 -7.315 ;
        RECT 242.595 -7.645 242.925 -7.315 ;
        RECT 241.235 -7.645 241.565 -7.315 ;
        RECT 239.875 -7.645 240.205 -7.315 ;
        RECT 238.515 -7.645 238.845 -7.315 ;
        RECT 237.155 -7.645 237.485 -7.315 ;
        RECT 235.795 -7.645 236.125 -7.315 ;
        RECT 234.435 -7.645 234.765 -7.315 ;
        RECT 233.075 -7.645 233.405 -7.315 ;
        RECT 231.715 -7.645 232.045 -7.315 ;
        RECT 230.355 -7.645 230.685 -7.315 ;
        RECT 228.995 -7.645 229.325 -7.315 ;
        RECT 227.635 -7.645 227.965 -7.315 ;
        RECT 226.275 -7.645 226.605 -7.315 ;
        RECT 224.915 -7.645 225.245 -7.315 ;
        RECT 223.555 -7.645 223.885 -7.315 ;
        RECT 222.195 -7.645 222.525 -7.315 ;
        RECT 220.835 -7.645 221.165 -7.315 ;
        RECT 219.475 -7.645 219.805 -7.315 ;
        RECT 218.115 -7.645 218.445 -7.315 ;
        RECT 216.755 -7.645 217.085 -7.315 ;
        RECT 215.395 -7.645 215.725 -7.315 ;
        RECT 214.035 -7.645 214.365 -7.315 ;
        RECT 212.675 -7.645 213.005 -7.315 ;
        RECT 211.315 -7.645 211.645 -7.315 ;
        RECT 209.955 -7.645 210.285 -7.315 ;
        RECT 208.595 -7.645 208.925 -7.315 ;
        RECT 207.235 -7.645 207.565 -7.315 ;
        RECT 205.875 -7.645 206.205 -7.315 ;
        RECT 204.515 -7.645 204.845 -7.315 ;
        RECT 203.155 -7.645 203.485 -7.315 ;
        RECT 201.795 -7.645 202.125 -7.315 ;
        RECT 200.435 -7.645 200.765 -7.315 ;
        RECT 199.075 -7.645 199.405 -7.315 ;
        RECT 197.715 -7.645 198.045 -7.315 ;
        RECT 196.355 -7.645 196.685 -7.315 ;
        RECT 194.995 -7.645 195.325 -7.315 ;
        RECT 193.635 -7.645 193.965 -7.315 ;
        RECT 192.275 -7.645 192.605 -7.315 ;
        RECT 190.915 -7.645 191.245 -7.315 ;
        RECT 189.555 -7.645 189.885 -7.315 ;
        RECT 188.195 -7.645 188.525 -7.315 ;
        RECT 186.835 -7.645 187.165 -7.315 ;
        RECT 185.475 -7.645 185.805 -7.315 ;
        RECT 184.115 -7.645 184.445 -7.315 ;
        RECT 182.755 -7.645 183.085 -7.315 ;
        RECT 181.395 -7.645 181.725 -7.315 ;
        RECT 180.035 -7.645 180.365 -7.315 ;
        RECT 178.675 -7.645 179.005 -7.315 ;
        RECT 177.315 -7.645 177.645 -7.315 ;
        RECT 175.955 -7.645 176.285 -7.315 ;
        RECT 174.595 -7.645 174.925 -7.315 ;
        RECT 173.235 -7.645 173.565 -7.315 ;
        RECT 171.875 -7.645 172.205 -7.315 ;
        RECT 170.515 -7.645 170.845 -7.315 ;
        RECT 169.155 -7.645 169.485 -7.315 ;
        RECT 167.795 -7.645 168.125 -7.315 ;
        RECT 166.435 -7.645 166.765 -7.315 ;
        RECT 165.075 -7.645 165.405 -7.315 ;
        RECT 163.715 -7.645 164.045 -7.315 ;
        RECT 162.355 -7.645 162.685 -7.315 ;
        RECT 160.995 -7.645 161.325 -7.315 ;
        RECT 159.635 -7.645 159.965 -7.315 ;
        RECT 158.275 -7.645 158.605 -7.315 ;
        RECT 156.915 -7.645 157.245 -7.315 ;
        RECT 155.555 -7.645 155.885 -7.315 ;
        RECT 154.195 -7.645 154.525 -7.315 ;
        RECT 152.835 -7.645 153.165 -7.315 ;
        RECT 151.475 -7.645 151.805 -7.315 ;
        RECT 150.115 -7.645 150.445 -7.315 ;
        RECT 148.755 -7.645 149.085 -7.315 ;
        RECT 147.395 -7.645 147.725 -7.315 ;
        RECT 146.035 -7.645 146.365 -7.315 ;
        RECT 144.675 -7.645 145.005 -7.315 ;
        RECT 143.315 -7.645 143.645 -7.315 ;
        RECT 141.955 -7.645 142.285 -7.315 ;
        RECT 140.595 -7.645 140.925 -7.315 ;
        RECT 139.235 -7.645 139.565 -7.315 ;
        RECT 137.875 -7.645 138.205 -7.315 ;
        RECT 136.515 -7.645 136.845 -7.315 ;
        RECT 135.155 -7.645 135.485 -7.315 ;
        RECT 133.795 -7.645 134.125 -7.315 ;
        RECT 132.435 -7.645 132.765 -7.315 ;
        RECT 131.075 -7.645 131.405 -7.315 ;
        RECT 129.715 -7.645 130.045 -7.315 ;
        RECT 128.355 -7.645 128.685 -7.315 ;
        RECT 126.995 -7.645 127.325 -7.315 ;
        RECT 125.635 -7.645 125.965 -7.315 ;
        RECT 124.275 -7.645 124.605 -7.315 ;
        RECT 122.915 -7.645 123.245 -7.315 ;
        RECT 121.555 -7.645 121.885 -7.315 ;
        RECT 120.195 -7.645 120.525 -7.315 ;
        RECT 118.835 -7.645 119.165 -7.315 ;
        RECT 117.475 -7.645 117.805 -7.315 ;
        RECT 116.115 -7.645 116.445 -7.315 ;
        RECT 114.755 -7.645 115.085 -7.315 ;
        RECT 113.395 -7.645 113.725 -7.315 ;
        RECT 112.035 -7.645 112.365 -7.315 ;
        RECT 110.675 -7.645 111.005 -7.315 ;
        RECT 109.315 -7.645 109.645 -7.315 ;
        RECT 107.955 -7.645 108.285 -7.315 ;
        RECT 106.595 -7.645 106.925 -7.315 ;
        RECT 105.235 -7.645 105.565 -7.315 ;
        RECT 103.875 -7.645 104.205 -7.315 ;
        RECT 102.515 -7.645 102.845 -7.315 ;
        RECT 101.155 -7.645 101.485 -7.315 ;
        RECT 99.795 -7.645 100.125 -7.315 ;
        RECT 98.435 -7.645 98.765 -7.315 ;
        RECT 97.075 -7.645 97.405 -7.315 ;
        RECT 95.715 -7.645 96.045 -7.315 ;
        RECT 94.355 -7.645 94.685 -7.315 ;
        RECT 92.995 -7.645 93.325 -7.315 ;
        RECT 91.635 -7.645 91.965 -7.315 ;
        RECT 90.275 -7.645 90.605 -7.315 ;
        RECT 88.915 -7.645 89.245 -7.315 ;
        RECT 87.555 -7.645 87.885 -7.315 ;
        RECT 86.195 -7.645 86.525 -7.315 ;
        RECT 84.835 -7.645 85.165 -7.315 ;
        RECT 83.475 -7.645 83.805 -7.315 ;
        RECT 82.115 -7.645 82.445 -7.315 ;
        RECT 80.755 -7.645 81.085 -7.315 ;
        RECT 79.395 -7.645 79.725 -7.315 ;
        RECT 78.035 -7.645 78.365 -7.315 ;
        RECT 76.675 -7.645 77.005 -7.315 ;
        RECT 75.315 -7.645 75.645 -7.315 ;
        RECT 73.955 -7.645 74.285 -7.315 ;
        RECT 72.595 -7.645 72.925 -7.315 ;
        RECT 71.235 -7.645 71.565 -7.315 ;
        RECT 69.875 -7.645 70.205 -7.315 ;
        RECT 68.515 -7.645 68.845 -7.315 ;
        RECT 67.155 -7.645 67.485 -7.315 ;
        RECT 65.795 -7.645 66.125 -7.315 ;
        RECT 64.435 -7.645 64.765 -7.315 ;
        RECT 63.075 -7.645 63.405 -7.315 ;
        RECT 61.715 -7.645 62.045 -7.315 ;
        RECT 60.355 -7.645 60.685 -7.315 ;
        RECT 58.995 -7.645 59.325 -7.315 ;
        RECT 57.635 -7.645 57.965 -7.315 ;
        RECT 56.275 -7.645 56.605 -7.315 ;
        RECT 54.915 -7.645 55.245 -7.315 ;
        RECT 53.555 -7.645 53.885 -7.315 ;
        RECT 52.195 -7.645 52.525 -7.315 ;
        RECT 50.835 -7.645 51.165 -7.315 ;
        RECT 49.475 -7.645 49.805 -7.315 ;
        RECT 48.115 -7.645 48.445 -7.315 ;
        RECT 46.755 -7.645 47.085 -7.315 ;
        RECT 45.395 -7.645 45.725 -7.315 ;
        RECT 44.035 -7.645 44.365 -7.315 ;
        RECT 42.675 -7.645 43.005 -7.315 ;
        RECT 41.315 -7.645 41.645 -7.315 ;
        RECT 39.955 -7.645 40.285 -7.315 ;
        RECT 38.595 -7.645 38.925 -7.315 ;
        RECT 37.235 -7.645 37.565 -7.315 ;
        RECT 35.875 -7.645 36.205 -7.315 ;
        RECT 34.515 -7.645 34.845 -7.315 ;
        RECT 33.155 -7.645 33.485 -7.315 ;
        RECT 31.795 -7.645 32.125 -7.315 ;
        RECT 30.435 -7.645 30.765 -7.315 ;
        RECT 29.075 -7.645 29.405 -7.315 ;
        RECT 27.715 -7.645 28.045 -7.315 ;
        RECT 26.355 -7.645 26.685 -7.315 ;
        RECT 24.995 -7.645 25.325 -7.315 ;
        RECT 23.635 -7.645 23.965 -7.315 ;
        RECT 22.275 -7.645 22.605 -7.315 ;
        RECT 20.915 -7.645 21.245 -7.315 ;
        RECT 19.555 -7.645 19.885 -7.315 ;
        RECT 18.195 -7.645 18.525 -7.315 ;
        RECT 16.835 -7.645 17.165 -7.315 ;
        RECT 15.475 -7.645 15.805 -7.315 ;
        RECT 14.115 -7.645 14.445 -7.315 ;
        RECT 12.755 -7.645 13.085 -7.315 ;
        RECT 11.395 -7.645 11.725 -7.315 ;
        RECT 10.035 -7.645 10.365 -7.315 ;
        RECT 8.675 -7.645 9.005 -7.315 ;
        RECT 7.315 -7.645 7.645 -7.315 ;
        RECT 5.955 -7.645 6.285 -7.315 ;
        RECT 4.595 -7.645 4.925 -7.315 ;
        RECT 3.235 -7.645 3.565 -7.315 ;
        RECT 1.875 -7.645 2.205 -7.315 ;
        RECT 0.515 -7.645 0.845 -7.315 ;
        RECT -0.845 -7.645 -0.515 -7.315 ;
        RECT 678.125 -7.64 954.88 -7.32 ;
        RECT 953.875 -7.645 954.205 -7.315 ;
        RECT 952.515 -7.645 952.845 -7.315 ;
        RECT 951.155 -7.645 951.485 -7.315 ;
        RECT 949.795 -7.645 950.125 -7.315 ;
        RECT 948.435 -7.645 948.765 -7.315 ;
        RECT 947.075 -7.645 947.405 -7.315 ;
        RECT 945.715 -7.645 946.045 -7.315 ;
        RECT 944.355 -7.645 944.685 -7.315 ;
        RECT 942.995 -7.645 943.325 -7.315 ;
        RECT 941.635 -7.645 941.965 -7.315 ;
        RECT 940.275 -7.645 940.605 -7.315 ;
        RECT 938.915 -7.645 939.245 -7.315 ;
        RECT 937.555 -7.645 937.885 -7.315 ;
        RECT 936.195 -7.645 936.525 -7.315 ;
        RECT 934.835 -7.645 935.165 -7.315 ;
        RECT 933.475 -7.645 933.805 -7.315 ;
        RECT 932.115 -7.645 932.445 -7.315 ;
        RECT 930.755 -7.645 931.085 -7.315 ;
        RECT 929.395 -7.645 929.725 -7.315 ;
        RECT 928.035 -7.645 928.365 -7.315 ;
        RECT 926.675 -7.645 927.005 -7.315 ;
        RECT 925.315 -7.645 925.645 -7.315 ;
        RECT 923.955 -7.645 924.285 -7.315 ;
        RECT 922.595 -7.645 922.925 -7.315 ;
        RECT 921.235 -7.645 921.565 -7.315 ;
        RECT 919.875 -7.645 920.205 -7.315 ;
        RECT 918.515 -7.645 918.845 -7.315 ;
        RECT 917.155 -7.645 917.485 -7.315 ;
        RECT 915.795 -7.645 916.125 -7.315 ;
        RECT 914.435 -7.645 914.765 -7.315 ;
        RECT 913.075 -7.645 913.405 -7.315 ;
        RECT 911.715 -7.645 912.045 -7.315 ;
        RECT 910.355 -7.645 910.685 -7.315 ;
        RECT 908.995 -7.645 909.325 -7.315 ;
        RECT 907.635 -7.645 907.965 -7.315 ;
        RECT 906.275 -7.645 906.605 -7.315 ;
        RECT 904.915 -7.645 905.245 -7.315 ;
        RECT 903.555 -7.645 903.885 -7.315 ;
        RECT 902.195 -7.645 902.525 -7.315 ;
        RECT 900.835 -7.645 901.165 -7.315 ;
        RECT 899.475 -7.645 899.805 -7.315 ;
        RECT 898.115 -7.645 898.445 -7.315 ;
        RECT 896.755 -7.645 897.085 -7.315 ;
        RECT 895.395 -7.645 895.725 -7.315 ;
        RECT 894.035 -7.645 894.365 -7.315 ;
        RECT 892.675 -7.645 893.005 -7.315 ;
        RECT 891.315 -7.645 891.645 -7.315 ;
        RECT 889.955 -7.645 890.285 -7.315 ;
        RECT 888.595 -7.645 888.925 -7.315 ;
        RECT 887.235 -7.645 887.565 -7.315 ;
        RECT 885.875 -7.645 886.205 -7.315 ;
        RECT 884.515 -7.645 884.845 -7.315 ;
        RECT 883.155 -7.645 883.485 -7.315 ;
        RECT 881.795 -7.645 882.125 -7.315 ;
        RECT 880.435 -7.645 880.765 -7.315 ;
        RECT 879.075 -7.645 879.405 -7.315 ;
        RECT 877.715 -7.645 878.045 -7.315 ;
        RECT 876.355 -7.645 876.685 -7.315 ;
        RECT 874.995 -7.645 875.325 -7.315 ;
        RECT 873.635 -7.645 873.965 -7.315 ;
        RECT 872.275 -7.645 872.605 -7.315 ;
        RECT 870.915 -7.645 871.245 -7.315 ;
        RECT 869.555 -7.645 869.885 -7.315 ;
        RECT 868.195 -7.645 868.525 -7.315 ;
        RECT 866.835 -7.645 867.165 -7.315 ;
        RECT 865.475 -7.645 865.805 -7.315 ;
        RECT 864.115 -7.645 864.445 -7.315 ;
        RECT 862.755 -7.645 863.085 -7.315 ;
        RECT 861.395 -7.645 861.725 -7.315 ;
        RECT 860.035 -7.645 860.365 -7.315 ;
        RECT 858.675 -7.645 859.005 -7.315 ;
        RECT 857.315 -7.645 857.645 -7.315 ;
        RECT 855.955 -7.645 856.285 -7.315 ;
        RECT 854.595 -7.645 854.925 -7.315 ;
        RECT 853.235 -7.645 853.565 -7.315 ;
        RECT 851.875 -7.645 852.205 -7.315 ;
        RECT 850.515 -7.645 850.845 -7.315 ;
        RECT 849.155 -7.645 849.485 -7.315 ;
        RECT 847.795 -7.645 848.125 -7.315 ;
        RECT 846.435 -7.645 846.765 -7.315 ;
        RECT 845.075 -7.645 845.405 -7.315 ;
        RECT 843.715 -7.645 844.045 -7.315 ;
        RECT 842.355 -7.645 842.685 -7.315 ;
        RECT 840.995 -7.645 841.325 -7.315 ;
        RECT 839.635 -7.645 839.965 -7.315 ;
        RECT 838.275 -7.645 838.605 -7.315 ;
        RECT 836.915 -7.645 837.245 -7.315 ;
        RECT 835.555 -7.645 835.885 -7.315 ;
        RECT 834.195 -7.645 834.525 -7.315 ;
        RECT 832.835 -7.645 833.165 -7.315 ;
        RECT 831.475 -7.645 831.805 -7.315 ;
        RECT 830.115 -7.645 830.445 -7.315 ;
        RECT 828.755 -7.645 829.085 -7.315 ;
        RECT 827.395 -7.645 827.725 -7.315 ;
        RECT 826.035 -7.645 826.365 -7.315 ;
        RECT 824.675 -7.645 825.005 -7.315 ;
        RECT 823.315 -7.645 823.645 -7.315 ;
        RECT 821.955 -7.645 822.285 -7.315 ;
        RECT 820.595 -7.645 820.925 -7.315 ;
        RECT 819.235 -7.645 819.565 -7.315 ;
        RECT 817.875 -7.645 818.205 -7.315 ;
        RECT 816.515 -7.645 816.845 -7.315 ;
        RECT 815.155 -7.645 815.485 -7.315 ;
        RECT 813.795 -7.645 814.125 -7.315 ;
        RECT 812.435 -7.645 812.765 -7.315 ;
        RECT 811.075 -7.645 811.405 -7.315 ;
        RECT 809.715 -7.645 810.045 -7.315 ;
        RECT 808.355 -7.645 808.685 -7.315 ;
        RECT 806.995 -7.645 807.325 -7.315 ;
        RECT 805.635 -7.645 805.965 -7.315 ;
        RECT 804.275 -7.645 804.605 -7.315 ;
        RECT 802.915 -7.645 803.245 -7.315 ;
        RECT 801.555 -7.645 801.885 -7.315 ;
        RECT 800.195 -7.645 800.525 -7.315 ;
        RECT 798.835 -7.645 799.165 -7.315 ;
        RECT 797.475 -7.645 797.805 -7.315 ;
        RECT 796.115 -7.645 796.445 -7.315 ;
        RECT 794.755 -7.645 795.085 -7.315 ;
        RECT 793.395 -7.645 793.725 -7.315 ;
        RECT 792.035 -7.645 792.365 -7.315 ;
        RECT 790.675 -7.645 791.005 -7.315 ;
        RECT 789.315 -7.645 789.645 -7.315 ;
        RECT 787.955 -7.645 788.285 -7.315 ;
        RECT 786.595 -7.645 786.925 -7.315 ;
        RECT 785.235 -7.645 785.565 -7.315 ;
        RECT 783.875 -7.645 784.205 -7.315 ;
        RECT 782.515 -7.645 782.845 -7.315 ;
        RECT 781.155 -7.645 781.485 -7.315 ;
        RECT 779.795 -7.645 780.125 -7.315 ;
        RECT 778.435 -7.645 778.765 -7.315 ;
        RECT 777.075 -7.645 777.405 -7.315 ;
        RECT 775.715 -7.645 776.045 -7.315 ;
        RECT 774.355 -7.645 774.685 -7.315 ;
        RECT 772.995 -7.645 773.325 -7.315 ;
        RECT 771.635 -7.645 771.965 -7.315 ;
        RECT 770.275 -7.645 770.605 -7.315 ;
        RECT 768.915 -7.645 769.245 -7.315 ;
        RECT 767.555 -7.645 767.885 -7.315 ;
        RECT 766.195 -7.645 766.525 -7.315 ;
        RECT 764.835 -7.645 765.165 -7.315 ;
        RECT 763.475 -7.645 763.805 -7.315 ;
        RECT 762.115 -7.645 762.445 -7.315 ;
        RECT 760.755 -7.645 761.085 -7.315 ;
        RECT 759.395 -7.645 759.725 -7.315 ;
        RECT 758.035 -7.645 758.365 -7.315 ;
        RECT 756.675 -7.645 757.005 -7.315 ;
        RECT 755.315 -7.645 755.645 -7.315 ;
        RECT 753.955 -7.645 754.285 -7.315 ;
        RECT 752.595 -7.645 752.925 -7.315 ;
        RECT 751.235 -7.645 751.565 -7.315 ;
        RECT 749.875 -7.645 750.205 -7.315 ;
        RECT 748.515 -7.645 748.845 -7.315 ;
        RECT 747.155 -7.645 747.485 -7.315 ;
        RECT 745.795 -7.645 746.125 -7.315 ;
        RECT 744.435 -7.645 744.765 -7.315 ;
        RECT 743.075 -7.645 743.405 -7.315 ;
        RECT 741.715 -7.645 742.045 -7.315 ;
        RECT 740.355 -7.645 740.685 -7.315 ;
        RECT 738.995 -7.645 739.325 -7.315 ;
        RECT 737.635 -7.645 737.965 -7.315 ;
        RECT 736.275 -7.645 736.605 -7.315 ;
        RECT 734.915 -7.645 735.245 -7.315 ;
        RECT 733.555 -7.645 733.885 -7.315 ;
        RECT 732.195 -7.645 732.525 -7.315 ;
        RECT 730.835 -7.645 731.165 -7.315 ;
        RECT 729.475 -7.645 729.805 -7.315 ;
        RECT 728.115 -7.645 728.445 -7.315 ;
        RECT 726.755 -7.645 727.085 -7.315 ;
        RECT 725.395 -7.645 725.725 -7.315 ;
        RECT 724.035 -7.645 724.365 -7.315 ;
        RECT 722.675 -7.645 723.005 -7.315 ;
        RECT 721.315 -7.645 721.645 -7.315 ;
        RECT 719.955 -7.645 720.285 -7.315 ;
        RECT 718.595 -7.645 718.925 -7.315 ;
        RECT 717.235 -7.645 717.565 -7.315 ;
        RECT 715.875 -7.645 716.205 -7.315 ;
        RECT 714.515 -7.645 714.845 -7.315 ;
        RECT 713.155 -7.645 713.485 -7.315 ;
        RECT 711.795 -7.645 712.125 -7.315 ;
        RECT 710.435 -7.645 710.765 -7.315 ;
        RECT 709.075 -7.645 709.405 -7.315 ;
        RECT 707.715 -7.645 708.045 -7.315 ;
        RECT 706.355 -7.645 706.685 -7.315 ;
        RECT 704.995 -7.645 705.325 -7.315 ;
        RECT 703.635 -7.645 703.965 -7.315 ;
        RECT 702.275 -7.645 702.605 -7.315 ;
        RECT 700.915 -7.645 701.245 -7.315 ;
        RECT 699.555 -7.645 699.885 -7.315 ;
        RECT 698.195 -7.645 698.525 -7.315 ;
        RECT 696.835 -7.645 697.165 -7.315 ;
        RECT 695.475 -7.645 695.805 -7.315 ;
        RECT 694.115 -7.645 694.445 -7.315 ;
        RECT 692.755 -7.645 693.085 -7.315 ;
        RECT 691.395 -7.645 691.725 -7.315 ;
        RECT 690.035 -7.645 690.365 -7.315 ;
        RECT 688.675 -7.645 689.005 -7.315 ;
        RECT 687.315 -7.645 687.645 -7.315 ;
        RECT 685.955 -7.645 686.285 -7.315 ;
        RECT 684.595 -7.645 684.925 -7.315 ;
        RECT 683.235 -7.645 683.565 -7.315 ;
        RECT 681.875 -7.645 682.205 -7.315 ;
        RECT 680.515 -7.645 680.845 -7.315 ;
        RECT 679.155 -7.645 679.485 -7.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -9.005 131.405 -8.675 ;
        RECT 129.715 -9.005 130.045 -8.675 ;
        RECT 128.355 -9.005 128.685 -8.675 ;
        RECT 126.995 -9.005 127.325 -8.675 ;
        RECT 125.635 -9.005 125.965 -8.675 ;
        RECT 124.275 -9.005 124.605 -8.675 ;
        RECT 122.915 -9.005 123.245 -8.675 ;
        RECT 121.555 -9.005 121.885 -8.675 ;
        RECT 120.195 -9.005 120.525 -8.675 ;
        RECT 118.835 -9.005 119.165 -8.675 ;
        RECT 117.475 -9.005 117.805 -8.675 ;
        RECT 116.115 -9.005 116.445 -8.675 ;
        RECT 114.755 -9.005 115.085 -8.675 ;
        RECT 113.395 -9.005 113.725 -8.675 ;
        RECT 112.035 -9.005 112.365 -8.675 ;
        RECT 110.675 -9.005 111.005 -8.675 ;
        RECT 109.315 -9.005 109.645 -8.675 ;
        RECT 107.955 -9.005 108.285 -8.675 ;
        RECT 106.595 -9.005 106.925 -8.675 ;
        RECT 105.235 -9.005 105.565 -8.675 ;
        RECT 103.875 -9.005 104.205 -8.675 ;
        RECT 102.515 -9.005 102.845 -8.675 ;
        RECT 101.155 -9.005 101.485 -8.675 ;
        RECT 99.795 -9.005 100.125 -8.675 ;
        RECT 98.435 -9.005 98.765 -8.675 ;
        RECT 97.075 -9.005 97.405 -8.675 ;
        RECT 95.715 -9.005 96.045 -8.675 ;
        RECT 94.355 -9.005 94.685 -8.675 ;
        RECT 92.995 -9.005 93.325 -8.675 ;
        RECT 91.635 -9.005 91.965 -8.675 ;
        RECT 90.275 -9.005 90.605 -8.675 ;
        RECT 88.915 -9.005 89.245 -8.675 ;
        RECT 87.555 -9.005 87.885 -8.675 ;
        RECT 86.195 -9.005 86.525 -8.675 ;
        RECT 84.835 -9.005 85.165 -8.675 ;
        RECT 83.475 -9.005 83.805 -8.675 ;
        RECT 82.115 -9.005 82.445 -8.675 ;
        RECT 80.755 -9.005 81.085 -8.675 ;
        RECT 79.395 -9.005 79.725 -8.675 ;
        RECT 78.035 -9.005 78.365 -8.675 ;
        RECT 76.675 -9.005 77.005 -8.675 ;
        RECT 75.315 -9.005 75.645 -8.675 ;
        RECT 73.955 -9.005 74.285 -8.675 ;
        RECT 72.595 -9.005 72.925 -8.675 ;
        RECT 71.235 -9.005 71.565 -8.675 ;
        RECT 69.875 -9.005 70.205 -8.675 ;
        RECT 68.515 -9.005 68.845 -8.675 ;
        RECT 67.155 -9.005 67.485 -8.675 ;
        RECT 65.795 -9.005 66.125 -8.675 ;
        RECT 64.435 -9.005 64.765 -8.675 ;
        RECT 63.075 -9.005 63.405 -8.675 ;
        RECT 61.715 -9.005 62.045 -8.675 ;
        RECT 60.355 -9.005 60.685 -8.675 ;
        RECT 58.995 -9.005 59.325 -8.675 ;
        RECT 57.635 -9.005 57.965 -8.675 ;
        RECT 56.275 -9.005 56.605 -8.675 ;
        RECT 54.915 -9.005 55.245 -8.675 ;
        RECT 53.555 -9.005 53.885 -8.675 ;
        RECT 52.195 -9.005 52.525 -8.675 ;
        RECT 50.835 -9.005 51.165 -8.675 ;
        RECT 49.475 -9.005 49.805 -8.675 ;
        RECT 48.115 -9.005 48.445 -8.675 ;
        RECT 46.755 -9.005 47.085 -8.675 ;
        RECT 45.395 -9.005 45.725 -8.675 ;
        RECT 44.035 -9.005 44.365 -8.675 ;
        RECT 42.675 -9.005 43.005 -8.675 ;
        RECT 41.315 -9.005 41.645 -8.675 ;
        RECT 39.955 -9.005 40.285 -8.675 ;
        RECT 38.595 -9.005 38.925 -8.675 ;
        RECT 37.235 -9.005 37.565 -8.675 ;
        RECT 35.875 -9.005 36.205 -8.675 ;
        RECT 34.515 -9.005 34.845 -8.675 ;
        RECT 33.155 -9.005 33.485 -8.675 ;
        RECT 31.795 -9.005 32.125 -8.675 ;
        RECT 30.435 -9.005 30.765 -8.675 ;
        RECT 29.075 -9.005 29.405 -8.675 ;
        RECT 27.715 -9.005 28.045 -8.675 ;
        RECT 26.355 -9.005 26.685 -8.675 ;
        RECT 24.995 -9.005 25.325 -8.675 ;
        RECT 23.635 -9.005 23.965 -8.675 ;
        RECT 22.275 -9.005 22.605 -8.675 ;
        RECT 20.915 -9.005 21.245 -8.675 ;
        RECT 19.555 -9.005 19.885 -8.675 ;
        RECT 18.195 -9.005 18.525 -8.675 ;
        RECT 16.835 -9.005 17.165 -8.675 ;
        RECT 15.475 -9.005 15.805 -8.675 ;
        RECT 14.115 -9.005 14.445 -8.675 ;
        RECT 12.755 -9.005 13.085 -8.675 ;
        RECT 11.395 -9.005 11.725 -8.675 ;
        RECT 10.035 -9.005 10.365 -8.675 ;
        RECT 8.675 -9.005 9.005 -8.675 ;
        RECT 7.315 -9.005 7.645 -8.675 ;
        RECT 5.955 -9.005 6.285 -8.675 ;
        RECT 4.595 -9.005 4.925 -8.675 ;
        RECT 3.235 -9.005 3.565 -8.675 ;
        RECT 1.875 -9.005 2.205 -8.675 ;
        RECT 0.515 -9.005 0.845 -8.675 ;
        RECT -0.845 -9.005 -0.515 -8.675 ;
        RECT 677.795 -9.005 678.125 -8.675 ;
        RECT -1.52 -9 678.125 -8.68 ;
        RECT 676.435 -9.005 676.765 -8.675 ;
        RECT 675.075 -9.005 675.405 -8.675 ;
        RECT 673.715 -9.005 674.045 -8.675 ;
        RECT 672.355 -9.005 672.685 -8.675 ;
        RECT 670.995 -9.005 671.325 -8.675 ;
        RECT 669.635 -9.005 669.965 -8.675 ;
        RECT 668.275 -9.005 668.605 -8.675 ;
        RECT 666.915 -9.005 667.245 -8.675 ;
        RECT 665.555 -9.005 665.885 -8.675 ;
        RECT 664.195 -9.005 664.525 -8.675 ;
        RECT 662.835 -9.005 663.165 -8.675 ;
        RECT 661.475 -9.005 661.805 -8.675 ;
        RECT 660.115 -9.005 660.445 -8.675 ;
        RECT 658.755 -9.005 659.085 -8.675 ;
        RECT 657.395 -9.005 657.725 -8.675 ;
        RECT 656.035 -9.005 656.365 -8.675 ;
        RECT 654.675 -9.005 655.005 -8.675 ;
        RECT 653.315 -9.005 653.645 -8.675 ;
        RECT 651.955 -9.005 652.285 -8.675 ;
        RECT 650.595 -9.005 650.925 -8.675 ;
        RECT 649.235 -9.005 649.565 -8.675 ;
        RECT 647.875 -9.005 648.205 -8.675 ;
        RECT 646.515 -9.005 646.845 -8.675 ;
        RECT 645.155 -9.005 645.485 -8.675 ;
        RECT 643.795 -9.005 644.125 -8.675 ;
        RECT 642.435 -9.005 642.765 -8.675 ;
        RECT 641.075 -9.005 641.405 -8.675 ;
        RECT 639.715 -9.005 640.045 -8.675 ;
        RECT 638.355 -9.005 638.685 -8.675 ;
        RECT 636.995 -9.005 637.325 -8.675 ;
        RECT 635.635 -9.005 635.965 -8.675 ;
        RECT 634.275 -9.005 634.605 -8.675 ;
        RECT 632.915 -9.005 633.245 -8.675 ;
        RECT 631.555 -9.005 631.885 -8.675 ;
        RECT 630.195 -9.005 630.525 -8.675 ;
        RECT 628.835 -9.005 629.165 -8.675 ;
        RECT 627.475 -9.005 627.805 -8.675 ;
        RECT 626.115 -9.005 626.445 -8.675 ;
        RECT 624.755 -9.005 625.085 -8.675 ;
        RECT 623.395 -9.005 623.725 -8.675 ;
        RECT 622.035 -9.005 622.365 -8.675 ;
        RECT 620.675 -9.005 621.005 -8.675 ;
        RECT 619.315 -9.005 619.645 -8.675 ;
        RECT 617.955 -9.005 618.285 -8.675 ;
        RECT 616.595 -9.005 616.925 -8.675 ;
        RECT 615.235 -9.005 615.565 -8.675 ;
        RECT 613.875 -9.005 614.205 -8.675 ;
        RECT 612.515 -9.005 612.845 -8.675 ;
        RECT 611.155 -9.005 611.485 -8.675 ;
        RECT 609.795 -9.005 610.125 -8.675 ;
        RECT 608.435 -9.005 608.765 -8.675 ;
        RECT 607.075 -9.005 607.405 -8.675 ;
        RECT 605.715 -9.005 606.045 -8.675 ;
        RECT 604.355 -9.005 604.685 -8.675 ;
        RECT 602.995 -9.005 603.325 -8.675 ;
        RECT 601.635 -9.005 601.965 -8.675 ;
        RECT 600.275 -9.005 600.605 -8.675 ;
        RECT 598.915 -9.005 599.245 -8.675 ;
        RECT 597.555 -9.005 597.885 -8.675 ;
        RECT 596.195 -9.005 596.525 -8.675 ;
        RECT 594.835 -9.005 595.165 -8.675 ;
        RECT 593.475 -9.005 593.805 -8.675 ;
        RECT 592.115 -9.005 592.445 -8.675 ;
        RECT 590.755 -9.005 591.085 -8.675 ;
        RECT 589.395 -9.005 589.725 -8.675 ;
        RECT 588.035 -9.005 588.365 -8.675 ;
        RECT 586.675 -9.005 587.005 -8.675 ;
        RECT 585.315 -9.005 585.645 -8.675 ;
        RECT 583.955 -9.005 584.285 -8.675 ;
        RECT 582.595 -9.005 582.925 -8.675 ;
        RECT 581.235 -9.005 581.565 -8.675 ;
        RECT 579.875 -9.005 580.205 -8.675 ;
        RECT 578.515 -9.005 578.845 -8.675 ;
        RECT 577.155 -9.005 577.485 -8.675 ;
        RECT 575.795 -9.005 576.125 -8.675 ;
        RECT 574.435 -9.005 574.765 -8.675 ;
        RECT 573.075 -9.005 573.405 -8.675 ;
        RECT 571.715 -9.005 572.045 -8.675 ;
        RECT 570.355 -9.005 570.685 -8.675 ;
        RECT 568.995 -9.005 569.325 -8.675 ;
        RECT 567.635 -9.005 567.965 -8.675 ;
        RECT 566.275 -9.005 566.605 -8.675 ;
        RECT 564.915 -9.005 565.245 -8.675 ;
        RECT 563.555 -9.005 563.885 -8.675 ;
        RECT 562.195 -9.005 562.525 -8.675 ;
        RECT 560.835 -9.005 561.165 -8.675 ;
        RECT 559.475 -9.005 559.805 -8.675 ;
        RECT 558.115 -9.005 558.445 -8.675 ;
        RECT 556.755 -9.005 557.085 -8.675 ;
        RECT 555.395 -9.005 555.725 -8.675 ;
        RECT 554.035 -9.005 554.365 -8.675 ;
        RECT 552.675 -9.005 553.005 -8.675 ;
        RECT 551.315 -9.005 551.645 -8.675 ;
        RECT 549.955 -9.005 550.285 -8.675 ;
        RECT 548.595 -9.005 548.925 -8.675 ;
        RECT 547.235 -9.005 547.565 -8.675 ;
        RECT 545.875 -9.005 546.205 -8.675 ;
        RECT 544.515 -9.005 544.845 -8.675 ;
        RECT 543.155 -9.005 543.485 -8.675 ;
        RECT 541.795 -9.005 542.125 -8.675 ;
        RECT 540.435 -9.005 540.765 -8.675 ;
        RECT 539.075 -9.005 539.405 -8.675 ;
        RECT 537.715 -9.005 538.045 -8.675 ;
        RECT 536.355 -9.005 536.685 -8.675 ;
        RECT 534.995 -9.005 535.325 -8.675 ;
        RECT 533.635 -9.005 533.965 -8.675 ;
        RECT 532.275 -9.005 532.605 -8.675 ;
        RECT 530.915 -9.005 531.245 -8.675 ;
        RECT 529.555 -9.005 529.885 -8.675 ;
        RECT 528.195 -9.005 528.525 -8.675 ;
        RECT 526.835 -9.005 527.165 -8.675 ;
        RECT 525.475 -9.005 525.805 -8.675 ;
        RECT 524.115 -9.005 524.445 -8.675 ;
        RECT 522.755 -9.005 523.085 -8.675 ;
        RECT 521.395 -9.005 521.725 -8.675 ;
        RECT 520.035 -9.005 520.365 -8.675 ;
        RECT 518.675 -9.005 519.005 -8.675 ;
        RECT 517.315 -9.005 517.645 -8.675 ;
        RECT 515.955 -9.005 516.285 -8.675 ;
        RECT 514.595 -9.005 514.925 -8.675 ;
        RECT 513.235 -9.005 513.565 -8.675 ;
        RECT 511.875 -9.005 512.205 -8.675 ;
        RECT 510.515 -9.005 510.845 -8.675 ;
        RECT 509.155 -9.005 509.485 -8.675 ;
        RECT 507.795 -9.005 508.125 -8.675 ;
        RECT 506.435 -9.005 506.765 -8.675 ;
        RECT 505.075 -9.005 505.405 -8.675 ;
        RECT 503.715 -9.005 504.045 -8.675 ;
        RECT 502.355 -9.005 502.685 -8.675 ;
        RECT 500.995 -9.005 501.325 -8.675 ;
        RECT 499.635 -9.005 499.965 -8.675 ;
        RECT 498.275 -9.005 498.605 -8.675 ;
        RECT 496.915 -9.005 497.245 -8.675 ;
        RECT 495.555 -9.005 495.885 -8.675 ;
        RECT 494.195 -9.005 494.525 -8.675 ;
        RECT 492.835 -9.005 493.165 -8.675 ;
        RECT 491.475 -9.005 491.805 -8.675 ;
        RECT 490.115 -9.005 490.445 -8.675 ;
        RECT 488.755 -9.005 489.085 -8.675 ;
        RECT 487.395 -9.005 487.725 -8.675 ;
        RECT 486.035 -9.005 486.365 -8.675 ;
        RECT 484.675 -9.005 485.005 -8.675 ;
        RECT 483.315 -9.005 483.645 -8.675 ;
        RECT 481.955 -9.005 482.285 -8.675 ;
        RECT 480.595 -9.005 480.925 -8.675 ;
        RECT 479.235 -9.005 479.565 -8.675 ;
        RECT 477.875 -9.005 478.205 -8.675 ;
        RECT 476.515 -9.005 476.845 -8.675 ;
        RECT 475.155 -9.005 475.485 -8.675 ;
        RECT 473.795 -9.005 474.125 -8.675 ;
        RECT 472.435 -9.005 472.765 -8.675 ;
        RECT 471.075 -9.005 471.405 -8.675 ;
        RECT 469.715 -9.005 470.045 -8.675 ;
        RECT 468.355 -9.005 468.685 -8.675 ;
        RECT 466.995 -9.005 467.325 -8.675 ;
        RECT 465.635 -9.005 465.965 -8.675 ;
        RECT 464.275 -9.005 464.605 -8.675 ;
        RECT 462.915 -9.005 463.245 -8.675 ;
        RECT 461.555 -9.005 461.885 -8.675 ;
        RECT 460.195 -9.005 460.525 -8.675 ;
        RECT 458.835 -9.005 459.165 -8.675 ;
        RECT 457.475 -9.005 457.805 -8.675 ;
        RECT 456.115 -9.005 456.445 -8.675 ;
        RECT 454.755 -9.005 455.085 -8.675 ;
        RECT 453.395 -9.005 453.725 -8.675 ;
        RECT 452.035 -9.005 452.365 -8.675 ;
        RECT 450.675 -9.005 451.005 -8.675 ;
        RECT 449.315 -9.005 449.645 -8.675 ;
        RECT 447.955 -9.005 448.285 -8.675 ;
        RECT 446.595 -9.005 446.925 -8.675 ;
        RECT 445.235 -9.005 445.565 -8.675 ;
        RECT 443.875 -9.005 444.205 -8.675 ;
        RECT 442.515 -9.005 442.845 -8.675 ;
        RECT 441.155 -9.005 441.485 -8.675 ;
        RECT 439.795 -9.005 440.125 -8.675 ;
        RECT 438.435 -9.005 438.765 -8.675 ;
        RECT 437.075 -9.005 437.405 -8.675 ;
        RECT 435.715 -9.005 436.045 -8.675 ;
        RECT 434.355 -9.005 434.685 -8.675 ;
        RECT 432.995 -9.005 433.325 -8.675 ;
        RECT 431.635 -9.005 431.965 -8.675 ;
        RECT 430.275 -9.005 430.605 -8.675 ;
        RECT 428.915 -9.005 429.245 -8.675 ;
        RECT 427.555 -9.005 427.885 -8.675 ;
        RECT 426.195 -9.005 426.525 -8.675 ;
        RECT 424.835 -9.005 425.165 -8.675 ;
        RECT 423.475 -9.005 423.805 -8.675 ;
        RECT 422.115 -9.005 422.445 -8.675 ;
        RECT 420.755 -9.005 421.085 -8.675 ;
        RECT 419.395 -9.005 419.725 -8.675 ;
        RECT 418.035 -9.005 418.365 -8.675 ;
        RECT 416.675 -9.005 417.005 -8.675 ;
        RECT 415.315 -9.005 415.645 -8.675 ;
        RECT 413.955 -9.005 414.285 -8.675 ;
        RECT 412.595 -9.005 412.925 -8.675 ;
        RECT 411.235 -9.005 411.565 -8.675 ;
        RECT 409.875 -9.005 410.205 -8.675 ;
        RECT 408.515 -9.005 408.845 -8.675 ;
        RECT 407.155 -9.005 407.485 -8.675 ;
        RECT 405.795 -9.005 406.125 -8.675 ;
        RECT 404.435 -9.005 404.765 -8.675 ;
        RECT 403.075 -9.005 403.405 -8.675 ;
        RECT 401.715 -9.005 402.045 -8.675 ;
        RECT 400.355 -9.005 400.685 -8.675 ;
        RECT 398.995 -9.005 399.325 -8.675 ;
        RECT 397.635 -9.005 397.965 -8.675 ;
        RECT 396.275 -9.005 396.605 -8.675 ;
        RECT 394.915 -9.005 395.245 -8.675 ;
        RECT 393.555 -9.005 393.885 -8.675 ;
        RECT 392.195 -9.005 392.525 -8.675 ;
        RECT 390.835 -9.005 391.165 -8.675 ;
        RECT 389.475 -9.005 389.805 -8.675 ;
        RECT 388.115 -9.005 388.445 -8.675 ;
        RECT 386.755 -9.005 387.085 -8.675 ;
        RECT 385.395 -9.005 385.725 -8.675 ;
        RECT 384.035 -9.005 384.365 -8.675 ;
        RECT 382.675 -9.005 383.005 -8.675 ;
        RECT 381.315 -9.005 381.645 -8.675 ;
        RECT 379.955 -9.005 380.285 -8.675 ;
        RECT 378.595 -9.005 378.925 -8.675 ;
        RECT 377.235 -9.005 377.565 -8.675 ;
        RECT 375.875 -9.005 376.205 -8.675 ;
        RECT 374.515 -9.005 374.845 -8.675 ;
        RECT 373.155 -9.005 373.485 -8.675 ;
        RECT 371.795 -9.005 372.125 -8.675 ;
        RECT 370.435 -9.005 370.765 -8.675 ;
        RECT 369.075 -9.005 369.405 -8.675 ;
        RECT 367.715 -9.005 368.045 -8.675 ;
        RECT 366.355 -9.005 366.685 -8.675 ;
        RECT 364.995 -9.005 365.325 -8.675 ;
        RECT 363.635 -9.005 363.965 -8.675 ;
        RECT 362.275 -9.005 362.605 -8.675 ;
        RECT 360.915 -9.005 361.245 -8.675 ;
        RECT 359.555 -9.005 359.885 -8.675 ;
        RECT 358.195 -9.005 358.525 -8.675 ;
        RECT 356.835 -9.005 357.165 -8.675 ;
        RECT 355.475 -9.005 355.805 -8.675 ;
        RECT 354.115 -9.005 354.445 -8.675 ;
        RECT 352.755 -9.005 353.085 -8.675 ;
        RECT 351.395 -9.005 351.725 -8.675 ;
        RECT 350.035 -9.005 350.365 -8.675 ;
        RECT 348.675 -9.005 349.005 -8.675 ;
        RECT 347.315 -9.005 347.645 -8.675 ;
        RECT 345.955 -9.005 346.285 -8.675 ;
        RECT 344.595 -9.005 344.925 -8.675 ;
        RECT 343.235 -9.005 343.565 -8.675 ;
        RECT 341.875 -9.005 342.205 -8.675 ;
        RECT 340.515 -9.005 340.845 -8.675 ;
        RECT 339.155 -9.005 339.485 -8.675 ;
        RECT 337.795 -9.005 338.125 -8.675 ;
        RECT 336.435 -9.005 336.765 -8.675 ;
        RECT 335.075 -9.005 335.405 -8.675 ;
        RECT 333.715 -9.005 334.045 -8.675 ;
        RECT 332.355 -9.005 332.685 -8.675 ;
        RECT 330.995 -9.005 331.325 -8.675 ;
        RECT 329.635 -9.005 329.965 -8.675 ;
        RECT 328.275 -9.005 328.605 -8.675 ;
        RECT 326.915 -9.005 327.245 -8.675 ;
        RECT 325.555 -9.005 325.885 -8.675 ;
        RECT 324.195 -9.005 324.525 -8.675 ;
        RECT 322.835 -9.005 323.165 -8.675 ;
        RECT 321.475 -9.005 321.805 -8.675 ;
        RECT 320.115 -9.005 320.445 -8.675 ;
        RECT 318.755 -9.005 319.085 -8.675 ;
        RECT 317.395 -9.005 317.725 -8.675 ;
        RECT 316.035 -9.005 316.365 -8.675 ;
        RECT 314.675 -9.005 315.005 -8.675 ;
        RECT 313.315 -9.005 313.645 -8.675 ;
        RECT 311.955 -9.005 312.285 -8.675 ;
        RECT 310.595 -9.005 310.925 -8.675 ;
        RECT 309.235 -9.005 309.565 -8.675 ;
        RECT 307.875 -9.005 308.205 -8.675 ;
        RECT 306.515 -9.005 306.845 -8.675 ;
        RECT 305.155 -9.005 305.485 -8.675 ;
        RECT 303.795 -9.005 304.125 -8.675 ;
        RECT 302.435 -9.005 302.765 -8.675 ;
        RECT 301.075 -9.005 301.405 -8.675 ;
        RECT 299.715 -9.005 300.045 -8.675 ;
        RECT 298.355 -9.005 298.685 -8.675 ;
        RECT 296.995 -9.005 297.325 -8.675 ;
        RECT 295.635 -9.005 295.965 -8.675 ;
        RECT 294.275 -9.005 294.605 -8.675 ;
        RECT 292.915 -9.005 293.245 -8.675 ;
        RECT 291.555 -9.005 291.885 -8.675 ;
        RECT 290.195 -9.005 290.525 -8.675 ;
        RECT 288.835 -9.005 289.165 -8.675 ;
        RECT 287.475 -9.005 287.805 -8.675 ;
        RECT 286.115 -9.005 286.445 -8.675 ;
        RECT 284.755 -9.005 285.085 -8.675 ;
        RECT 283.395 -9.005 283.725 -8.675 ;
        RECT 282.035 -9.005 282.365 -8.675 ;
        RECT 280.675 -9.005 281.005 -8.675 ;
        RECT 279.315 -9.005 279.645 -8.675 ;
        RECT 277.955 -9.005 278.285 -8.675 ;
        RECT 276.595 -9.005 276.925 -8.675 ;
        RECT 275.235 -9.005 275.565 -8.675 ;
        RECT 273.875 -9.005 274.205 -8.675 ;
        RECT 272.515 -9.005 272.845 -8.675 ;
        RECT 271.155 -9.005 271.485 -8.675 ;
        RECT 269.795 -9.005 270.125 -8.675 ;
        RECT 268.435 -9.005 268.765 -8.675 ;
        RECT 267.075 -9.005 267.405 -8.675 ;
        RECT 265.715 -9.005 266.045 -8.675 ;
        RECT 264.355 -9.005 264.685 -8.675 ;
        RECT 262.995 -9.005 263.325 -8.675 ;
        RECT 261.635 -9.005 261.965 -8.675 ;
        RECT 260.275 -9.005 260.605 -8.675 ;
        RECT 258.915 -9.005 259.245 -8.675 ;
        RECT 257.555 -9.005 257.885 -8.675 ;
        RECT 256.195 -9.005 256.525 -8.675 ;
        RECT 254.835 -9.005 255.165 -8.675 ;
        RECT 253.475 -9.005 253.805 -8.675 ;
        RECT 252.115 -9.005 252.445 -8.675 ;
        RECT 250.755 -9.005 251.085 -8.675 ;
        RECT 249.395 -9.005 249.725 -8.675 ;
        RECT 248.035 -9.005 248.365 -8.675 ;
        RECT 246.675 -9.005 247.005 -8.675 ;
        RECT 245.315 -9.005 245.645 -8.675 ;
        RECT 243.955 -9.005 244.285 -8.675 ;
        RECT 242.595 -9.005 242.925 -8.675 ;
        RECT 241.235 -9.005 241.565 -8.675 ;
        RECT 239.875 -9.005 240.205 -8.675 ;
        RECT 238.515 -9.005 238.845 -8.675 ;
        RECT 237.155 -9.005 237.485 -8.675 ;
        RECT 235.795 -9.005 236.125 -8.675 ;
        RECT 234.435 -9.005 234.765 -8.675 ;
        RECT 233.075 -9.005 233.405 -8.675 ;
        RECT 231.715 -9.005 232.045 -8.675 ;
        RECT 230.355 -9.005 230.685 -8.675 ;
        RECT 228.995 -9.005 229.325 -8.675 ;
        RECT 227.635 -9.005 227.965 -8.675 ;
        RECT 226.275 -9.005 226.605 -8.675 ;
        RECT 224.915 -9.005 225.245 -8.675 ;
        RECT 223.555 -9.005 223.885 -8.675 ;
        RECT 222.195 -9.005 222.525 -8.675 ;
        RECT 220.835 -9.005 221.165 -8.675 ;
        RECT 219.475 -9.005 219.805 -8.675 ;
        RECT 218.115 -9.005 218.445 -8.675 ;
        RECT 216.755 -9.005 217.085 -8.675 ;
        RECT 215.395 -9.005 215.725 -8.675 ;
        RECT 214.035 -9.005 214.365 -8.675 ;
        RECT 212.675 -9.005 213.005 -8.675 ;
        RECT 211.315 -9.005 211.645 -8.675 ;
        RECT 209.955 -9.005 210.285 -8.675 ;
        RECT 208.595 -9.005 208.925 -8.675 ;
        RECT 207.235 -9.005 207.565 -8.675 ;
        RECT 205.875 -9.005 206.205 -8.675 ;
        RECT 204.515 -9.005 204.845 -8.675 ;
        RECT 203.155 -9.005 203.485 -8.675 ;
        RECT 201.795 -9.005 202.125 -8.675 ;
        RECT 200.435 -9.005 200.765 -8.675 ;
        RECT 199.075 -9.005 199.405 -8.675 ;
        RECT 197.715 -9.005 198.045 -8.675 ;
        RECT 196.355 -9.005 196.685 -8.675 ;
        RECT 194.995 -9.005 195.325 -8.675 ;
        RECT 193.635 -9.005 193.965 -8.675 ;
        RECT 192.275 -9.005 192.605 -8.675 ;
        RECT 190.915 -9.005 191.245 -8.675 ;
        RECT 189.555 -9.005 189.885 -8.675 ;
        RECT 188.195 -9.005 188.525 -8.675 ;
        RECT 186.835 -9.005 187.165 -8.675 ;
        RECT 185.475 -9.005 185.805 -8.675 ;
        RECT 184.115 -9.005 184.445 -8.675 ;
        RECT 182.755 -9.005 183.085 -8.675 ;
        RECT 181.395 -9.005 181.725 -8.675 ;
        RECT 180.035 -9.005 180.365 -8.675 ;
        RECT 178.675 -9.005 179.005 -8.675 ;
        RECT 177.315 -9.005 177.645 -8.675 ;
        RECT 175.955 -9.005 176.285 -8.675 ;
        RECT 174.595 -9.005 174.925 -8.675 ;
        RECT 173.235 -9.005 173.565 -8.675 ;
        RECT 171.875 -9.005 172.205 -8.675 ;
        RECT 170.515 -9.005 170.845 -8.675 ;
        RECT 169.155 -9.005 169.485 -8.675 ;
        RECT 167.795 -9.005 168.125 -8.675 ;
        RECT 166.435 -9.005 166.765 -8.675 ;
        RECT 165.075 -9.005 165.405 -8.675 ;
        RECT 163.715 -9.005 164.045 -8.675 ;
        RECT 162.355 -9.005 162.685 -8.675 ;
        RECT 160.995 -9.005 161.325 -8.675 ;
        RECT 159.635 -9.005 159.965 -8.675 ;
        RECT 158.275 -9.005 158.605 -8.675 ;
        RECT 156.915 -9.005 157.245 -8.675 ;
        RECT 155.555 -9.005 155.885 -8.675 ;
        RECT 154.195 -9.005 154.525 -8.675 ;
        RECT 152.835 -9.005 153.165 -8.675 ;
        RECT 151.475 -9.005 151.805 -8.675 ;
        RECT 150.115 -9.005 150.445 -8.675 ;
        RECT 148.755 -9.005 149.085 -8.675 ;
        RECT 147.395 -9.005 147.725 -8.675 ;
        RECT 146.035 -9.005 146.365 -8.675 ;
        RECT 144.675 -9.005 145.005 -8.675 ;
        RECT 143.315 -9.005 143.645 -8.675 ;
        RECT 141.955 -9.005 142.285 -8.675 ;
        RECT 140.595 -9.005 140.925 -8.675 ;
        RECT 139.235 -9.005 139.565 -8.675 ;
        RECT 137.875 -9.005 138.205 -8.675 ;
        RECT 136.515 -9.005 136.845 -8.675 ;
        RECT 135.155 -9.005 135.485 -8.675 ;
        RECT 133.795 -9.005 134.125 -8.675 ;
        RECT 132.435 -9.005 132.765 -8.675 ;
        RECT 678.125 -9 954.88 -8.68 ;
        RECT 953.875 -9.005 954.205 -8.675 ;
        RECT 952.515 -9.005 952.845 -8.675 ;
        RECT 951.155 -9.005 951.485 -8.675 ;
        RECT 949.795 -9.005 950.125 -8.675 ;
        RECT 948.435 -9.005 948.765 -8.675 ;
        RECT 947.075 -9.005 947.405 -8.675 ;
        RECT 945.715 -9.005 946.045 -8.675 ;
        RECT 944.355 -9.005 944.685 -8.675 ;
        RECT 942.995 -9.005 943.325 -8.675 ;
        RECT 941.635 -9.005 941.965 -8.675 ;
        RECT 940.275 -9.005 940.605 -8.675 ;
        RECT 938.915 -9.005 939.245 -8.675 ;
        RECT 937.555 -9.005 937.885 -8.675 ;
        RECT 936.195 -9.005 936.525 -8.675 ;
        RECT 934.835 -9.005 935.165 -8.675 ;
        RECT 933.475 -9.005 933.805 -8.675 ;
        RECT 932.115 -9.005 932.445 -8.675 ;
        RECT 930.755 -9.005 931.085 -8.675 ;
        RECT 929.395 -9.005 929.725 -8.675 ;
        RECT 928.035 -9.005 928.365 -8.675 ;
        RECT 926.675 -9.005 927.005 -8.675 ;
        RECT 925.315 -9.005 925.645 -8.675 ;
        RECT 923.955 -9.005 924.285 -8.675 ;
        RECT 922.595 -9.005 922.925 -8.675 ;
        RECT 921.235 -9.005 921.565 -8.675 ;
        RECT 919.875 -9.005 920.205 -8.675 ;
        RECT 918.515 -9.005 918.845 -8.675 ;
        RECT 917.155 -9.005 917.485 -8.675 ;
        RECT 915.795 -9.005 916.125 -8.675 ;
        RECT 914.435 -9.005 914.765 -8.675 ;
        RECT 913.075 -9.005 913.405 -8.675 ;
        RECT 911.715 -9.005 912.045 -8.675 ;
        RECT 910.355 -9.005 910.685 -8.675 ;
        RECT 908.995 -9.005 909.325 -8.675 ;
        RECT 907.635 -9.005 907.965 -8.675 ;
        RECT 906.275 -9.005 906.605 -8.675 ;
        RECT 904.915 -9.005 905.245 -8.675 ;
        RECT 903.555 -9.005 903.885 -8.675 ;
        RECT 902.195 -9.005 902.525 -8.675 ;
        RECT 900.835 -9.005 901.165 -8.675 ;
        RECT 899.475 -9.005 899.805 -8.675 ;
        RECT 898.115 -9.005 898.445 -8.675 ;
        RECT 896.755 -9.005 897.085 -8.675 ;
        RECT 895.395 -9.005 895.725 -8.675 ;
        RECT 894.035 -9.005 894.365 -8.675 ;
        RECT 892.675 -9.005 893.005 -8.675 ;
        RECT 891.315 -9.005 891.645 -8.675 ;
        RECT 889.955 -9.005 890.285 -8.675 ;
        RECT 888.595 -9.005 888.925 -8.675 ;
        RECT 887.235 -9.005 887.565 -8.675 ;
        RECT 885.875 -9.005 886.205 -8.675 ;
        RECT 884.515 -9.005 884.845 -8.675 ;
        RECT 883.155 -9.005 883.485 -8.675 ;
        RECT 881.795 -9.005 882.125 -8.675 ;
        RECT 880.435 -9.005 880.765 -8.675 ;
        RECT 879.075 -9.005 879.405 -8.675 ;
        RECT 877.715 -9.005 878.045 -8.675 ;
        RECT 876.355 -9.005 876.685 -8.675 ;
        RECT 874.995 -9.005 875.325 -8.675 ;
        RECT 873.635 -9.005 873.965 -8.675 ;
        RECT 872.275 -9.005 872.605 -8.675 ;
        RECT 870.915 -9.005 871.245 -8.675 ;
        RECT 869.555 -9.005 869.885 -8.675 ;
        RECT 868.195 -9.005 868.525 -8.675 ;
        RECT 866.835 -9.005 867.165 -8.675 ;
        RECT 865.475 -9.005 865.805 -8.675 ;
        RECT 864.115 -9.005 864.445 -8.675 ;
        RECT 862.755 -9.005 863.085 -8.675 ;
        RECT 861.395 -9.005 861.725 -8.675 ;
        RECT 860.035 -9.005 860.365 -8.675 ;
        RECT 858.675 -9.005 859.005 -8.675 ;
        RECT 857.315 -9.005 857.645 -8.675 ;
        RECT 855.955 -9.005 856.285 -8.675 ;
        RECT 854.595 -9.005 854.925 -8.675 ;
        RECT 853.235 -9.005 853.565 -8.675 ;
        RECT 851.875 -9.005 852.205 -8.675 ;
        RECT 850.515 -9.005 850.845 -8.675 ;
        RECT 849.155 -9.005 849.485 -8.675 ;
        RECT 847.795 -9.005 848.125 -8.675 ;
        RECT 846.435 -9.005 846.765 -8.675 ;
        RECT 845.075 -9.005 845.405 -8.675 ;
        RECT 843.715 -9.005 844.045 -8.675 ;
        RECT 842.355 -9.005 842.685 -8.675 ;
        RECT 840.995 -9.005 841.325 -8.675 ;
        RECT 839.635 -9.005 839.965 -8.675 ;
        RECT 838.275 -9.005 838.605 -8.675 ;
        RECT 836.915 -9.005 837.245 -8.675 ;
        RECT 835.555 -9.005 835.885 -8.675 ;
        RECT 834.195 -9.005 834.525 -8.675 ;
        RECT 832.835 -9.005 833.165 -8.675 ;
        RECT 831.475 -9.005 831.805 -8.675 ;
        RECT 830.115 -9.005 830.445 -8.675 ;
        RECT 828.755 -9.005 829.085 -8.675 ;
        RECT 827.395 -9.005 827.725 -8.675 ;
        RECT 826.035 -9.005 826.365 -8.675 ;
        RECT 824.675 -9.005 825.005 -8.675 ;
        RECT 823.315 -9.005 823.645 -8.675 ;
        RECT 821.955 -9.005 822.285 -8.675 ;
        RECT 820.595 -9.005 820.925 -8.675 ;
        RECT 819.235 -9.005 819.565 -8.675 ;
        RECT 817.875 -9.005 818.205 -8.675 ;
        RECT 816.515 -9.005 816.845 -8.675 ;
        RECT 815.155 -9.005 815.485 -8.675 ;
        RECT 813.795 -9.005 814.125 -8.675 ;
        RECT 812.435 -9.005 812.765 -8.675 ;
        RECT 811.075 -9.005 811.405 -8.675 ;
        RECT 809.715 -9.005 810.045 -8.675 ;
        RECT 808.355 -9.005 808.685 -8.675 ;
        RECT 806.995 -9.005 807.325 -8.675 ;
        RECT 805.635 -9.005 805.965 -8.675 ;
        RECT 804.275 -9.005 804.605 -8.675 ;
        RECT 802.915 -9.005 803.245 -8.675 ;
        RECT 801.555 -9.005 801.885 -8.675 ;
        RECT 800.195 -9.005 800.525 -8.675 ;
        RECT 798.835 -9.005 799.165 -8.675 ;
        RECT 797.475 -9.005 797.805 -8.675 ;
        RECT 796.115 -9.005 796.445 -8.675 ;
        RECT 794.755 -9.005 795.085 -8.675 ;
        RECT 793.395 -9.005 793.725 -8.675 ;
        RECT 792.035 -9.005 792.365 -8.675 ;
        RECT 790.675 -9.005 791.005 -8.675 ;
        RECT 789.315 -9.005 789.645 -8.675 ;
        RECT 787.955 -9.005 788.285 -8.675 ;
        RECT 786.595 -9.005 786.925 -8.675 ;
        RECT 785.235 -9.005 785.565 -8.675 ;
        RECT 783.875 -9.005 784.205 -8.675 ;
        RECT 782.515 -9.005 782.845 -8.675 ;
        RECT 781.155 -9.005 781.485 -8.675 ;
        RECT 779.795 -9.005 780.125 -8.675 ;
        RECT 778.435 -9.005 778.765 -8.675 ;
        RECT 777.075 -9.005 777.405 -8.675 ;
        RECT 775.715 -9.005 776.045 -8.675 ;
        RECT 774.355 -9.005 774.685 -8.675 ;
        RECT 772.995 -9.005 773.325 -8.675 ;
        RECT 771.635 -9.005 771.965 -8.675 ;
        RECT 770.275 -9.005 770.605 -8.675 ;
        RECT 768.915 -9.005 769.245 -8.675 ;
        RECT 767.555 -9.005 767.885 -8.675 ;
        RECT 766.195 -9.005 766.525 -8.675 ;
        RECT 764.835 -9.005 765.165 -8.675 ;
        RECT 763.475 -9.005 763.805 -8.675 ;
        RECT 762.115 -9.005 762.445 -8.675 ;
        RECT 760.755 -9.005 761.085 -8.675 ;
        RECT 759.395 -9.005 759.725 -8.675 ;
        RECT 758.035 -9.005 758.365 -8.675 ;
        RECT 756.675 -9.005 757.005 -8.675 ;
        RECT 755.315 -9.005 755.645 -8.675 ;
        RECT 753.955 -9.005 754.285 -8.675 ;
        RECT 752.595 -9.005 752.925 -8.675 ;
        RECT 751.235 -9.005 751.565 -8.675 ;
        RECT 749.875 -9.005 750.205 -8.675 ;
        RECT 748.515 -9.005 748.845 -8.675 ;
        RECT 747.155 -9.005 747.485 -8.675 ;
        RECT 745.795 -9.005 746.125 -8.675 ;
        RECT 744.435 -9.005 744.765 -8.675 ;
        RECT 743.075 -9.005 743.405 -8.675 ;
        RECT 741.715 -9.005 742.045 -8.675 ;
        RECT 740.355 -9.005 740.685 -8.675 ;
        RECT 738.995 -9.005 739.325 -8.675 ;
        RECT 737.635 -9.005 737.965 -8.675 ;
        RECT 736.275 -9.005 736.605 -8.675 ;
        RECT 734.915 -9.005 735.245 -8.675 ;
        RECT 733.555 -9.005 733.885 -8.675 ;
        RECT 732.195 -9.005 732.525 -8.675 ;
        RECT 730.835 -9.005 731.165 -8.675 ;
        RECT 729.475 -9.005 729.805 -8.675 ;
        RECT 728.115 -9.005 728.445 -8.675 ;
        RECT 726.755 -9.005 727.085 -8.675 ;
        RECT 725.395 -9.005 725.725 -8.675 ;
        RECT 724.035 -9.005 724.365 -8.675 ;
        RECT 722.675 -9.005 723.005 -8.675 ;
        RECT 721.315 -9.005 721.645 -8.675 ;
        RECT 719.955 -9.005 720.285 -8.675 ;
        RECT 718.595 -9.005 718.925 -8.675 ;
        RECT 717.235 -9.005 717.565 -8.675 ;
        RECT 715.875 -9.005 716.205 -8.675 ;
        RECT 714.515 -9.005 714.845 -8.675 ;
        RECT 713.155 -9.005 713.485 -8.675 ;
        RECT 711.795 -9.005 712.125 -8.675 ;
        RECT 710.435 -9.005 710.765 -8.675 ;
        RECT 709.075 -9.005 709.405 -8.675 ;
        RECT 707.715 -9.005 708.045 -8.675 ;
        RECT 706.355 -9.005 706.685 -8.675 ;
        RECT 704.995 -9.005 705.325 -8.675 ;
        RECT 703.635 -9.005 703.965 -8.675 ;
        RECT 702.275 -9.005 702.605 -8.675 ;
        RECT 700.915 -9.005 701.245 -8.675 ;
        RECT 699.555 -9.005 699.885 -8.675 ;
        RECT 698.195 -9.005 698.525 -8.675 ;
        RECT 696.835 -9.005 697.165 -8.675 ;
        RECT 695.475 -9.005 695.805 -8.675 ;
        RECT 694.115 -9.005 694.445 -8.675 ;
        RECT 692.755 -9.005 693.085 -8.675 ;
        RECT 691.395 -9.005 691.725 -8.675 ;
        RECT 690.035 -9.005 690.365 -8.675 ;
        RECT 688.675 -9.005 689.005 -8.675 ;
        RECT 687.315 -9.005 687.645 -8.675 ;
        RECT 685.955 -9.005 686.285 -8.675 ;
        RECT 684.595 -9.005 684.925 -8.675 ;
        RECT 683.235 -9.005 683.565 -8.675 ;
        RECT 681.875 -9.005 682.205 -8.675 ;
        RECT 680.515 -9.005 680.845 -8.675 ;
        RECT 679.155 -9.005 679.485 -8.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 -4.925 678.125 -4.595 ;
        RECT -1.52 -4.92 678.125 -4.6 ;
        RECT 676.435 -4.925 676.765 -4.595 ;
        RECT 675.075 -4.925 675.405 -4.595 ;
        RECT 673.715 -4.925 674.045 -4.595 ;
        RECT 672.355 -4.925 672.685 -4.595 ;
        RECT 670.995 -4.925 671.325 -4.595 ;
        RECT 669.635 -4.925 669.965 -4.595 ;
        RECT 668.275 -4.925 668.605 -4.595 ;
        RECT 666.915 -4.925 667.245 -4.595 ;
        RECT 665.555 -4.925 665.885 -4.595 ;
        RECT 664.195 -4.925 664.525 -4.595 ;
        RECT 662.835 -4.925 663.165 -4.595 ;
        RECT 661.475 -4.925 661.805 -4.595 ;
        RECT 660.115 -4.925 660.445 -4.595 ;
        RECT 658.755 -4.925 659.085 -4.595 ;
        RECT 657.395 -4.925 657.725 -4.595 ;
        RECT 656.035 -4.925 656.365 -4.595 ;
        RECT 654.675 -4.925 655.005 -4.595 ;
        RECT 653.315 -4.925 653.645 -4.595 ;
        RECT 651.955 -4.925 652.285 -4.595 ;
        RECT 650.595 -4.925 650.925 -4.595 ;
        RECT 649.235 -4.925 649.565 -4.595 ;
        RECT 647.875 -4.925 648.205 -4.595 ;
        RECT 646.515 -4.925 646.845 -4.595 ;
        RECT 645.155 -4.925 645.485 -4.595 ;
        RECT 643.795 -4.925 644.125 -4.595 ;
        RECT 642.435 -4.925 642.765 -4.595 ;
        RECT 641.075 -4.925 641.405 -4.595 ;
        RECT 639.715 -4.925 640.045 -4.595 ;
        RECT 638.355 -4.925 638.685 -4.595 ;
        RECT 636.995 -4.925 637.325 -4.595 ;
        RECT 635.635 -4.925 635.965 -4.595 ;
        RECT 634.275 -4.925 634.605 -4.595 ;
        RECT 632.915 -4.925 633.245 -4.595 ;
        RECT 631.555 -4.925 631.885 -4.595 ;
        RECT 630.195 -4.925 630.525 -4.595 ;
        RECT 628.835 -4.925 629.165 -4.595 ;
        RECT 627.475 -4.925 627.805 -4.595 ;
        RECT 626.115 -4.925 626.445 -4.595 ;
        RECT 624.755 -4.925 625.085 -4.595 ;
        RECT 623.395 -4.925 623.725 -4.595 ;
        RECT 622.035 -4.925 622.365 -4.595 ;
        RECT 620.675 -4.925 621.005 -4.595 ;
        RECT 619.315 -4.925 619.645 -4.595 ;
        RECT 617.955 -4.925 618.285 -4.595 ;
        RECT 616.595 -4.925 616.925 -4.595 ;
        RECT 615.235 -4.925 615.565 -4.595 ;
        RECT 613.875 -4.925 614.205 -4.595 ;
        RECT 612.515 -4.925 612.845 -4.595 ;
        RECT 611.155 -4.925 611.485 -4.595 ;
        RECT 609.795 -4.925 610.125 -4.595 ;
        RECT 608.435 -4.925 608.765 -4.595 ;
        RECT 607.075 -4.925 607.405 -4.595 ;
        RECT 605.715 -4.925 606.045 -4.595 ;
        RECT 604.355 -4.925 604.685 -4.595 ;
        RECT 602.995 -4.925 603.325 -4.595 ;
        RECT 601.635 -4.925 601.965 -4.595 ;
        RECT 600.275 -4.925 600.605 -4.595 ;
        RECT 598.915 -4.925 599.245 -4.595 ;
        RECT 597.555 -4.925 597.885 -4.595 ;
        RECT 596.195 -4.925 596.525 -4.595 ;
        RECT 594.835 -4.925 595.165 -4.595 ;
        RECT 593.475 -4.925 593.805 -4.595 ;
        RECT 592.115 -4.925 592.445 -4.595 ;
        RECT 590.755 -4.925 591.085 -4.595 ;
        RECT 589.395 -4.925 589.725 -4.595 ;
        RECT 588.035 -4.925 588.365 -4.595 ;
        RECT 586.675 -4.925 587.005 -4.595 ;
        RECT 585.315 -4.925 585.645 -4.595 ;
        RECT 583.955 -4.925 584.285 -4.595 ;
        RECT 582.595 -4.925 582.925 -4.595 ;
        RECT 581.235 -4.925 581.565 -4.595 ;
        RECT 579.875 -4.925 580.205 -4.595 ;
        RECT 578.515 -4.925 578.845 -4.595 ;
        RECT 577.155 -4.925 577.485 -4.595 ;
        RECT 575.795 -4.925 576.125 -4.595 ;
        RECT 574.435 -4.925 574.765 -4.595 ;
        RECT 573.075 -4.925 573.405 -4.595 ;
        RECT 571.715 -4.925 572.045 -4.595 ;
        RECT 570.355 -4.925 570.685 -4.595 ;
        RECT 568.995 -4.925 569.325 -4.595 ;
        RECT 567.635 -4.925 567.965 -4.595 ;
        RECT 566.275 -4.925 566.605 -4.595 ;
        RECT 564.915 -4.925 565.245 -4.595 ;
        RECT 563.555 -4.925 563.885 -4.595 ;
        RECT 562.195 -4.925 562.525 -4.595 ;
        RECT 560.835 -4.925 561.165 -4.595 ;
        RECT 559.475 -4.925 559.805 -4.595 ;
        RECT 558.115 -4.925 558.445 -4.595 ;
        RECT 556.755 -4.925 557.085 -4.595 ;
        RECT 555.395 -4.925 555.725 -4.595 ;
        RECT 554.035 -4.925 554.365 -4.595 ;
        RECT 552.675 -4.925 553.005 -4.595 ;
        RECT 551.315 -4.925 551.645 -4.595 ;
        RECT 549.955 -4.925 550.285 -4.595 ;
        RECT 548.595 -4.925 548.925 -4.595 ;
        RECT 547.235 -4.925 547.565 -4.595 ;
        RECT 545.875 -4.925 546.205 -4.595 ;
        RECT 544.515 -4.925 544.845 -4.595 ;
        RECT 543.155 -4.925 543.485 -4.595 ;
        RECT 541.795 -4.925 542.125 -4.595 ;
        RECT 540.435 -4.925 540.765 -4.595 ;
        RECT 539.075 -4.925 539.405 -4.595 ;
        RECT 537.715 -4.925 538.045 -4.595 ;
        RECT 536.355 -4.925 536.685 -4.595 ;
        RECT 534.995 -4.925 535.325 -4.595 ;
        RECT 533.635 -4.925 533.965 -4.595 ;
        RECT 532.275 -4.925 532.605 -4.595 ;
        RECT 530.915 -4.925 531.245 -4.595 ;
        RECT 529.555 -4.925 529.885 -4.595 ;
        RECT 528.195 -4.925 528.525 -4.595 ;
        RECT 526.835 -4.925 527.165 -4.595 ;
        RECT 525.475 -4.925 525.805 -4.595 ;
        RECT 524.115 -4.925 524.445 -4.595 ;
        RECT 522.755 -4.925 523.085 -4.595 ;
        RECT 521.395 -4.925 521.725 -4.595 ;
        RECT 520.035 -4.925 520.365 -4.595 ;
        RECT 518.675 -4.925 519.005 -4.595 ;
        RECT 517.315 -4.925 517.645 -4.595 ;
        RECT 515.955 -4.925 516.285 -4.595 ;
        RECT 514.595 -4.925 514.925 -4.595 ;
        RECT 513.235 -4.925 513.565 -4.595 ;
        RECT 511.875 -4.925 512.205 -4.595 ;
        RECT 510.515 -4.925 510.845 -4.595 ;
        RECT 509.155 -4.925 509.485 -4.595 ;
        RECT 507.795 -4.925 508.125 -4.595 ;
        RECT 506.435 -4.925 506.765 -4.595 ;
        RECT 505.075 -4.925 505.405 -4.595 ;
        RECT 503.715 -4.925 504.045 -4.595 ;
        RECT 502.355 -4.925 502.685 -4.595 ;
        RECT 500.995 -4.925 501.325 -4.595 ;
        RECT 499.635 -4.925 499.965 -4.595 ;
        RECT 498.275 -4.925 498.605 -4.595 ;
        RECT 496.915 -4.925 497.245 -4.595 ;
        RECT 495.555 -4.925 495.885 -4.595 ;
        RECT 494.195 -4.925 494.525 -4.595 ;
        RECT 492.835 -4.925 493.165 -4.595 ;
        RECT 491.475 -4.925 491.805 -4.595 ;
        RECT 490.115 -4.925 490.445 -4.595 ;
        RECT 488.755 -4.925 489.085 -4.595 ;
        RECT 487.395 -4.925 487.725 -4.595 ;
        RECT 486.035 -4.925 486.365 -4.595 ;
        RECT 484.675 -4.925 485.005 -4.595 ;
        RECT 483.315 -4.925 483.645 -4.595 ;
        RECT 481.955 -4.925 482.285 -4.595 ;
        RECT 480.595 -4.925 480.925 -4.595 ;
        RECT 479.235 -4.925 479.565 -4.595 ;
        RECT 477.875 -4.925 478.205 -4.595 ;
        RECT 476.515 -4.925 476.845 -4.595 ;
        RECT 475.155 -4.925 475.485 -4.595 ;
        RECT 473.795 -4.925 474.125 -4.595 ;
        RECT 472.435 -4.925 472.765 -4.595 ;
        RECT 471.075 -4.925 471.405 -4.595 ;
        RECT 469.715 -4.925 470.045 -4.595 ;
        RECT 468.355 -4.925 468.685 -4.595 ;
        RECT 466.995 -4.925 467.325 -4.595 ;
        RECT 465.635 -4.925 465.965 -4.595 ;
        RECT 464.275 -4.925 464.605 -4.595 ;
        RECT 462.915 -4.925 463.245 -4.595 ;
        RECT 461.555 -4.925 461.885 -4.595 ;
        RECT 460.195 -4.925 460.525 -4.595 ;
        RECT 458.835 -4.925 459.165 -4.595 ;
        RECT 457.475 -4.925 457.805 -4.595 ;
        RECT 456.115 -4.925 456.445 -4.595 ;
        RECT 454.755 -4.925 455.085 -4.595 ;
        RECT 453.395 -4.925 453.725 -4.595 ;
        RECT 452.035 -4.925 452.365 -4.595 ;
        RECT 450.675 -4.925 451.005 -4.595 ;
        RECT 449.315 -4.925 449.645 -4.595 ;
        RECT 447.955 -4.925 448.285 -4.595 ;
        RECT 446.595 -4.925 446.925 -4.595 ;
        RECT 445.235 -4.925 445.565 -4.595 ;
        RECT 443.875 -4.925 444.205 -4.595 ;
        RECT 442.515 -4.925 442.845 -4.595 ;
        RECT 441.155 -4.925 441.485 -4.595 ;
        RECT 439.795 -4.925 440.125 -4.595 ;
        RECT 438.435 -4.925 438.765 -4.595 ;
        RECT 437.075 -4.925 437.405 -4.595 ;
        RECT 435.715 -4.925 436.045 -4.595 ;
        RECT 434.355 -4.925 434.685 -4.595 ;
        RECT 432.995 -4.925 433.325 -4.595 ;
        RECT 431.635 -4.925 431.965 -4.595 ;
        RECT 430.275 -4.925 430.605 -4.595 ;
        RECT 428.915 -4.925 429.245 -4.595 ;
        RECT 427.555 -4.925 427.885 -4.595 ;
        RECT 426.195 -4.925 426.525 -4.595 ;
        RECT 424.835 -4.925 425.165 -4.595 ;
        RECT 423.475 -4.925 423.805 -4.595 ;
        RECT 422.115 -4.925 422.445 -4.595 ;
        RECT 420.755 -4.925 421.085 -4.595 ;
        RECT 419.395 -4.925 419.725 -4.595 ;
        RECT 418.035 -4.925 418.365 -4.595 ;
        RECT 416.675 -4.925 417.005 -4.595 ;
        RECT 415.315 -4.925 415.645 -4.595 ;
        RECT 413.955 -4.925 414.285 -4.595 ;
        RECT 412.595 -4.925 412.925 -4.595 ;
        RECT 411.235 -4.925 411.565 -4.595 ;
        RECT 409.875 -4.925 410.205 -4.595 ;
        RECT 408.515 -4.925 408.845 -4.595 ;
        RECT 407.155 -4.925 407.485 -4.595 ;
        RECT 405.795 -4.925 406.125 -4.595 ;
        RECT 404.435 -4.925 404.765 -4.595 ;
        RECT 403.075 -4.925 403.405 -4.595 ;
        RECT 401.715 -4.925 402.045 -4.595 ;
        RECT 400.355 -4.925 400.685 -4.595 ;
        RECT 398.995 -4.925 399.325 -4.595 ;
        RECT 397.635 -4.925 397.965 -4.595 ;
        RECT 396.275 -4.925 396.605 -4.595 ;
        RECT 394.915 -4.925 395.245 -4.595 ;
        RECT 393.555 -4.925 393.885 -4.595 ;
        RECT 392.195 -4.925 392.525 -4.595 ;
        RECT 390.835 -4.925 391.165 -4.595 ;
        RECT 389.475 -4.925 389.805 -4.595 ;
        RECT 388.115 -4.925 388.445 -4.595 ;
        RECT 386.755 -4.925 387.085 -4.595 ;
        RECT 385.395 -4.925 385.725 -4.595 ;
        RECT 384.035 -4.925 384.365 -4.595 ;
        RECT 382.675 -4.925 383.005 -4.595 ;
        RECT 381.315 -4.925 381.645 -4.595 ;
        RECT 379.955 -4.925 380.285 -4.595 ;
        RECT 378.595 -4.925 378.925 -4.595 ;
        RECT 377.235 -4.925 377.565 -4.595 ;
        RECT 375.875 -4.925 376.205 -4.595 ;
        RECT 374.515 -4.925 374.845 -4.595 ;
        RECT 373.155 -4.925 373.485 -4.595 ;
        RECT 371.795 -4.925 372.125 -4.595 ;
        RECT 370.435 -4.925 370.765 -4.595 ;
        RECT 369.075 -4.925 369.405 -4.595 ;
        RECT 367.715 -4.925 368.045 -4.595 ;
        RECT 366.355 -4.925 366.685 -4.595 ;
        RECT 364.995 -4.925 365.325 -4.595 ;
        RECT 363.635 -4.925 363.965 -4.595 ;
        RECT 362.275 -4.925 362.605 -4.595 ;
        RECT 360.915 -4.925 361.245 -4.595 ;
        RECT 359.555 -4.925 359.885 -4.595 ;
        RECT 358.195 -4.925 358.525 -4.595 ;
        RECT 356.835 -4.925 357.165 -4.595 ;
        RECT 355.475 -4.925 355.805 -4.595 ;
        RECT 354.115 -4.925 354.445 -4.595 ;
        RECT 352.755 -4.925 353.085 -4.595 ;
        RECT 351.395 -4.925 351.725 -4.595 ;
        RECT 350.035 -4.925 350.365 -4.595 ;
        RECT 348.675 -4.925 349.005 -4.595 ;
        RECT 347.315 -4.925 347.645 -4.595 ;
        RECT 345.955 -4.925 346.285 -4.595 ;
        RECT 344.595 -4.925 344.925 -4.595 ;
        RECT 343.235 -4.925 343.565 -4.595 ;
        RECT 341.875 -4.925 342.205 -4.595 ;
        RECT 340.515 -4.925 340.845 -4.595 ;
        RECT 339.155 -4.925 339.485 -4.595 ;
        RECT 337.795 -4.925 338.125 -4.595 ;
        RECT 336.435 -4.925 336.765 -4.595 ;
        RECT 335.075 -4.925 335.405 -4.595 ;
        RECT 333.715 -4.925 334.045 -4.595 ;
        RECT 332.355 -4.925 332.685 -4.595 ;
        RECT 330.995 -4.925 331.325 -4.595 ;
        RECT 329.635 -4.925 329.965 -4.595 ;
        RECT 328.275 -4.925 328.605 -4.595 ;
        RECT 326.915 -4.925 327.245 -4.595 ;
        RECT 325.555 -4.925 325.885 -4.595 ;
        RECT 324.195 -4.925 324.525 -4.595 ;
        RECT 322.835 -4.925 323.165 -4.595 ;
        RECT 321.475 -4.925 321.805 -4.595 ;
        RECT 320.115 -4.925 320.445 -4.595 ;
        RECT 318.755 -4.925 319.085 -4.595 ;
        RECT 317.395 -4.925 317.725 -4.595 ;
        RECT 316.035 -4.925 316.365 -4.595 ;
        RECT 314.675 -4.925 315.005 -4.595 ;
        RECT 313.315 -4.925 313.645 -4.595 ;
        RECT 311.955 -4.925 312.285 -4.595 ;
        RECT 310.595 -4.925 310.925 -4.595 ;
        RECT 309.235 -4.925 309.565 -4.595 ;
        RECT 307.875 -4.925 308.205 -4.595 ;
        RECT 306.515 -4.925 306.845 -4.595 ;
        RECT 305.155 -4.925 305.485 -4.595 ;
        RECT 303.795 -4.925 304.125 -4.595 ;
        RECT 302.435 -4.925 302.765 -4.595 ;
        RECT 301.075 -4.925 301.405 -4.595 ;
        RECT 299.715 -4.925 300.045 -4.595 ;
        RECT 298.355 -4.925 298.685 -4.595 ;
        RECT 296.995 -4.925 297.325 -4.595 ;
        RECT 295.635 -4.925 295.965 -4.595 ;
        RECT 294.275 -4.925 294.605 -4.595 ;
        RECT 292.915 -4.925 293.245 -4.595 ;
        RECT 291.555 -4.925 291.885 -4.595 ;
        RECT 290.195 -4.925 290.525 -4.595 ;
        RECT 288.835 -4.925 289.165 -4.595 ;
        RECT 287.475 -4.925 287.805 -4.595 ;
        RECT 286.115 -4.925 286.445 -4.595 ;
        RECT 284.755 -4.925 285.085 -4.595 ;
        RECT 283.395 -4.925 283.725 -4.595 ;
        RECT 282.035 -4.925 282.365 -4.595 ;
        RECT 280.675 -4.925 281.005 -4.595 ;
        RECT 279.315 -4.925 279.645 -4.595 ;
        RECT 277.955 -4.925 278.285 -4.595 ;
        RECT 276.595 -4.925 276.925 -4.595 ;
        RECT 275.235 -4.925 275.565 -4.595 ;
        RECT 273.875 -4.925 274.205 -4.595 ;
        RECT 272.515 -4.925 272.845 -4.595 ;
        RECT 271.155 -4.925 271.485 -4.595 ;
        RECT 269.795 -4.925 270.125 -4.595 ;
        RECT 268.435 -4.925 268.765 -4.595 ;
        RECT 267.075 -4.925 267.405 -4.595 ;
        RECT 265.715 -4.925 266.045 -4.595 ;
        RECT 264.355 -4.925 264.685 -4.595 ;
        RECT 262.995 -4.925 263.325 -4.595 ;
        RECT 261.635 -4.925 261.965 -4.595 ;
        RECT 260.275 -4.925 260.605 -4.595 ;
        RECT 258.915 -4.925 259.245 -4.595 ;
        RECT 257.555 -4.925 257.885 -4.595 ;
        RECT 256.195 -4.925 256.525 -4.595 ;
        RECT 254.835 -4.925 255.165 -4.595 ;
        RECT 253.475 -4.925 253.805 -4.595 ;
        RECT 252.115 -4.925 252.445 -4.595 ;
        RECT 250.755 -4.925 251.085 -4.595 ;
        RECT 249.395 -4.925 249.725 -4.595 ;
        RECT 248.035 -4.925 248.365 -4.595 ;
        RECT 246.675 -4.925 247.005 -4.595 ;
        RECT 245.315 -4.925 245.645 -4.595 ;
        RECT 243.955 -4.925 244.285 -4.595 ;
        RECT 242.595 -4.925 242.925 -4.595 ;
        RECT 241.235 -4.925 241.565 -4.595 ;
        RECT 239.875 -4.925 240.205 -4.595 ;
        RECT 238.515 -4.925 238.845 -4.595 ;
        RECT 237.155 -4.925 237.485 -4.595 ;
        RECT 235.795 -4.925 236.125 -4.595 ;
        RECT 234.435 -4.925 234.765 -4.595 ;
        RECT 233.075 -4.925 233.405 -4.595 ;
        RECT 231.715 -4.925 232.045 -4.595 ;
        RECT 230.355 -4.925 230.685 -4.595 ;
        RECT 228.995 -4.925 229.325 -4.595 ;
        RECT 227.635 -4.925 227.965 -4.595 ;
        RECT 226.275 -4.925 226.605 -4.595 ;
        RECT 224.915 -4.925 225.245 -4.595 ;
        RECT 223.555 -4.925 223.885 -4.595 ;
        RECT 222.195 -4.925 222.525 -4.595 ;
        RECT 220.835 -4.925 221.165 -4.595 ;
        RECT 219.475 -4.925 219.805 -4.595 ;
        RECT 218.115 -4.925 218.445 -4.595 ;
        RECT 216.755 -4.925 217.085 -4.595 ;
        RECT 215.395 -4.925 215.725 -4.595 ;
        RECT 214.035 -4.925 214.365 -4.595 ;
        RECT 212.675 -4.925 213.005 -4.595 ;
        RECT 211.315 -4.925 211.645 -4.595 ;
        RECT 209.955 -4.925 210.285 -4.595 ;
        RECT 208.595 -4.925 208.925 -4.595 ;
        RECT 207.235 -4.925 207.565 -4.595 ;
        RECT 205.875 -4.925 206.205 -4.595 ;
        RECT 204.515 -4.925 204.845 -4.595 ;
        RECT 203.155 -4.925 203.485 -4.595 ;
        RECT 201.795 -4.925 202.125 -4.595 ;
        RECT 200.435 -4.925 200.765 -4.595 ;
        RECT 199.075 -4.925 199.405 -4.595 ;
        RECT 197.715 -4.925 198.045 -4.595 ;
        RECT 196.355 -4.925 196.685 -4.595 ;
        RECT 194.995 -4.925 195.325 -4.595 ;
        RECT 193.635 -4.925 193.965 -4.595 ;
        RECT 192.275 -4.925 192.605 -4.595 ;
        RECT 190.915 -4.925 191.245 -4.595 ;
        RECT 189.555 -4.925 189.885 -4.595 ;
        RECT 188.195 -4.925 188.525 -4.595 ;
        RECT 186.835 -4.925 187.165 -4.595 ;
        RECT 185.475 -4.925 185.805 -4.595 ;
        RECT 184.115 -4.925 184.445 -4.595 ;
        RECT 182.755 -4.925 183.085 -4.595 ;
        RECT 181.395 -4.925 181.725 -4.595 ;
        RECT 180.035 -4.925 180.365 -4.595 ;
        RECT 178.675 -4.925 179.005 -4.595 ;
        RECT 177.315 -4.925 177.645 -4.595 ;
        RECT 175.955 -4.925 176.285 -4.595 ;
        RECT 174.595 -4.925 174.925 -4.595 ;
        RECT 173.235 -4.925 173.565 -4.595 ;
        RECT 171.875 -4.925 172.205 -4.595 ;
        RECT 170.515 -4.925 170.845 -4.595 ;
        RECT 169.155 -4.925 169.485 -4.595 ;
        RECT 167.795 -4.925 168.125 -4.595 ;
        RECT 166.435 -4.925 166.765 -4.595 ;
        RECT 165.075 -4.925 165.405 -4.595 ;
        RECT 163.715 -4.925 164.045 -4.595 ;
        RECT 162.355 -4.925 162.685 -4.595 ;
        RECT 160.995 -4.925 161.325 -4.595 ;
        RECT 159.635 -4.925 159.965 -4.595 ;
        RECT 158.275 -4.925 158.605 -4.595 ;
        RECT 156.915 -4.925 157.245 -4.595 ;
        RECT 155.555 -4.925 155.885 -4.595 ;
        RECT 154.195 -4.925 154.525 -4.595 ;
        RECT 152.835 -4.925 153.165 -4.595 ;
        RECT 151.475 -4.925 151.805 -4.595 ;
        RECT 150.115 -4.925 150.445 -4.595 ;
        RECT 148.755 -4.925 149.085 -4.595 ;
        RECT 147.395 -4.925 147.725 -4.595 ;
        RECT 146.035 -4.925 146.365 -4.595 ;
        RECT 144.675 -4.925 145.005 -4.595 ;
        RECT 143.315 -4.925 143.645 -4.595 ;
        RECT 141.955 -4.925 142.285 -4.595 ;
        RECT 140.595 -4.925 140.925 -4.595 ;
        RECT 139.235 -4.925 139.565 -4.595 ;
        RECT 137.875 -4.925 138.205 -4.595 ;
        RECT 136.515 -4.925 136.845 -4.595 ;
        RECT 135.155 -4.925 135.485 -4.595 ;
        RECT 133.795 -4.925 134.125 -4.595 ;
        RECT 132.435 -4.925 132.765 -4.595 ;
        RECT 131.075 -4.925 131.405 -4.595 ;
        RECT 129.715 -4.925 130.045 -4.595 ;
        RECT 128.355 -4.925 128.685 -4.595 ;
        RECT 126.995 -4.925 127.325 -4.595 ;
        RECT 125.635 -4.925 125.965 -4.595 ;
        RECT 124.275 -4.925 124.605 -4.595 ;
        RECT 122.915 -4.925 123.245 -4.595 ;
        RECT 121.555 -4.925 121.885 -4.595 ;
        RECT 120.195 -4.925 120.525 -4.595 ;
        RECT 118.835 -4.925 119.165 -4.595 ;
        RECT 117.475 -4.925 117.805 -4.595 ;
        RECT 116.115 -4.925 116.445 -4.595 ;
        RECT 114.755 -4.925 115.085 -4.595 ;
        RECT 113.395 -4.925 113.725 -4.595 ;
        RECT 112.035 -4.925 112.365 -4.595 ;
        RECT 110.675 -4.925 111.005 -4.595 ;
        RECT 109.315 -4.925 109.645 -4.595 ;
        RECT 107.955 -4.925 108.285 -4.595 ;
        RECT 106.595 -4.925 106.925 -4.595 ;
        RECT 105.235 -4.925 105.565 -4.595 ;
        RECT 103.875 -4.925 104.205 -4.595 ;
        RECT 102.515 -4.925 102.845 -4.595 ;
        RECT 101.155 -4.925 101.485 -4.595 ;
        RECT 99.795 -4.925 100.125 -4.595 ;
        RECT 98.435 -4.925 98.765 -4.595 ;
        RECT 97.075 -4.925 97.405 -4.595 ;
        RECT 95.715 -4.925 96.045 -4.595 ;
        RECT 94.355 -4.925 94.685 -4.595 ;
        RECT 92.995 -4.925 93.325 -4.595 ;
        RECT 91.635 -4.925 91.965 -4.595 ;
        RECT 90.275 -4.925 90.605 -4.595 ;
        RECT 88.915 -4.925 89.245 -4.595 ;
        RECT 87.555 -4.925 87.885 -4.595 ;
        RECT 86.195 -4.925 86.525 -4.595 ;
        RECT 84.835 -4.925 85.165 -4.595 ;
        RECT 83.475 -4.925 83.805 -4.595 ;
        RECT 82.115 -4.925 82.445 -4.595 ;
        RECT 80.755 -4.925 81.085 -4.595 ;
        RECT 79.395 -4.925 79.725 -4.595 ;
        RECT 78.035 -4.925 78.365 -4.595 ;
        RECT 76.675 -4.925 77.005 -4.595 ;
        RECT 75.315 -4.925 75.645 -4.595 ;
        RECT 73.955 -4.925 74.285 -4.595 ;
        RECT 72.595 -4.925 72.925 -4.595 ;
        RECT 71.235 -4.925 71.565 -4.595 ;
        RECT 69.875 -4.925 70.205 -4.595 ;
        RECT 68.515 -4.925 68.845 -4.595 ;
        RECT 67.155 -4.925 67.485 -4.595 ;
        RECT 65.795 -4.925 66.125 -4.595 ;
        RECT 64.435 -4.925 64.765 -4.595 ;
        RECT 63.075 -4.925 63.405 -4.595 ;
        RECT 61.715 -4.925 62.045 -4.595 ;
        RECT 60.355 -4.925 60.685 -4.595 ;
        RECT 58.995 -4.925 59.325 -4.595 ;
        RECT 57.635 -4.925 57.965 -4.595 ;
        RECT 56.275 -4.925 56.605 -4.595 ;
        RECT 54.915 -4.925 55.245 -4.595 ;
        RECT 53.555 -4.925 53.885 -4.595 ;
        RECT 52.195 -4.925 52.525 -4.595 ;
        RECT 50.835 -4.925 51.165 -4.595 ;
        RECT 49.475 -4.925 49.805 -4.595 ;
        RECT 48.115 -4.925 48.445 -4.595 ;
        RECT 46.755 -4.925 47.085 -4.595 ;
        RECT 45.395 -4.925 45.725 -4.595 ;
        RECT 44.035 -4.925 44.365 -4.595 ;
        RECT 42.675 -4.925 43.005 -4.595 ;
        RECT 41.315 -4.925 41.645 -4.595 ;
        RECT 39.955 -4.925 40.285 -4.595 ;
        RECT 38.595 -4.925 38.925 -4.595 ;
        RECT 37.235 -4.925 37.565 -4.595 ;
        RECT 35.875 -4.925 36.205 -4.595 ;
        RECT 34.515 -4.925 34.845 -4.595 ;
        RECT 33.155 -4.925 33.485 -4.595 ;
        RECT 31.795 -4.925 32.125 -4.595 ;
        RECT 30.435 -4.925 30.765 -4.595 ;
        RECT 29.075 -4.925 29.405 -4.595 ;
        RECT 27.715 -4.925 28.045 -4.595 ;
        RECT 26.355 -4.925 26.685 -4.595 ;
        RECT 24.995 -4.925 25.325 -4.595 ;
        RECT 23.635 -4.925 23.965 -4.595 ;
        RECT 22.275 -4.925 22.605 -4.595 ;
        RECT 20.915 -4.925 21.245 -4.595 ;
        RECT 19.555 -4.925 19.885 -4.595 ;
        RECT 18.195 -4.925 18.525 -4.595 ;
        RECT 16.835 -4.925 17.165 -4.595 ;
        RECT 15.475 -4.925 15.805 -4.595 ;
        RECT 14.115 -4.925 14.445 -4.595 ;
        RECT 12.755 -4.925 13.085 -4.595 ;
        RECT 11.395 -4.925 11.725 -4.595 ;
        RECT 10.035 -4.925 10.365 -4.595 ;
        RECT 8.675 -4.925 9.005 -4.595 ;
        RECT 7.315 -4.925 7.645 -4.595 ;
        RECT 5.955 -4.925 6.285 -4.595 ;
        RECT 4.595 -4.925 4.925 -4.595 ;
        RECT 3.235 -4.925 3.565 -4.595 ;
        RECT 1.875 -4.925 2.205 -4.595 ;
        RECT 0.515 -4.925 0.845 -4.595 ;
        RECT -0.845 -4.925 -0.515 -4.595 ;
        RECT 762.115 -4.925 762.445 -4.595 ;
        RECT 760.755 -4.925 761.085 -4.595 ;
        RECT 759.395 -4.925 759.725 -4.595 ;
        RECT 758.035 -4.925 758.365 -4.595 ;
        RECT 756.675 -4.925 757.005 -4.595 ;
        RECT 755.315 -4.925 755.645 -4.595 ;
        RECT 753.955 -4.925 754.285 -4.595 ;
        RECT 752.595 -4.925 752.925 -4.595 ;
        RECT 751.235 -4.925 751.565 -4.595 ;
        RECT 749.875 -4.925 750.205 -4.595 ;
        RECT 748.515 -4.925 748.845 -4.595 ;
        RECT 747.155 -4.925 747.485 -4.595 ;
        RECT 745.795 -4.925 746.125 -4.595 ;
        RECT 744.435 -4.925 744.765 -4.595 ;
        RECT 743.075 -4.925 743.405 -4.595 ;
        RECT 741.715 -4.925 742.045 -4.595 ;
        RECT 740.355 -4.925 740.685 -4.595 ;
        RECT 738.995 -4.925 739.325 -4.595 ;
        RECT 737.635 -4.925 737.965 -4.595 ;
        RECT 736.275 -4.925 736.605 -4.595 ;
        RECT 734.915 -4.925 735.245 -4.595 ;
        RECT 733.555 -4.925 733.885 -4.595 ;
        RECT 732.195 -4.925 732.525 -4.595 ;
        RECT 730.835 -4.925 731.165 -4.595 ;
        RECT 729.475 -4.925 729.805 -4.595 ;
        RECT 728.115 -4.925 728.445 -4.595 ;
        RECT 726.755 -4.925 727.085 -4.595 ;
        RECT 725.395 -4.925 725.725 -4.595 ;
        RECT 724.035 -4.925 724.365 -4.595 ;
        RECT 722.675 -4.925 723.005 -4.595 ;
        RECT 721.315 -4.925 721.645 -4.595 ;
        RECT 719.955 -4.925 720.285 -4.595 ;
        RECT 718.595 -4.925 718.925 -4.595 ;
        RECT 717.235 -4.925 717.565 -4.595 ;
        RECT 715.875 -4.925 716.205 -4.595 ;
        RECT 714.515 -4.925 714.845 -4.595 ;
        RECT 713.155 -4.925 713.485 -4.595 ;
        RECT 711.795 -4.925 712.125 -4.595 ;
        RECT 710.435 -4.925 710.765 -4.595 ;
        RECT 709.075 -4.925 709.405 -4.595 ;
        RECT 707.715 -4.925 708.045 -4.595 ;
        RECT 706.355 -4.925 706.685 -4.595 ;
        RECT 704.995 -4.925 705.325 -4.595 ;
        RECT 703.635 -4.925 703.965 -4.595 ;
        RECT 702.275 -4.925 702.605 -4.595 ;
        RECT 700.915 -4.925 701.245 -4.595 ;
        RECT 699.555 -4.925 699.885 -4.595 ;
        RECT 698.195 -4.925 698.525 -4.595 ;
        RECT 696.835 -4.925 697.165 -4.595 ;
        RECT 695.475 -4.925 695.805 -4.595 ;
        RECT 694.115 -4.925 694.445 -4.595 ;
        RECT 692.755 -4.925 693.085 -4.595 ;
        RECT 691.395 -4.925 691.725 -4.595 ;
        RECT 690.035 -4.925 690.365 -4.595 ;
        RECT 688.675 -4.925 689.005 -4.595 ;
        RECT 687.315 -4.925 687.645 -4.595 ;
        RECT 685.955 -4.925 686.285 -4.595 ;
        RECT 684.595 -4.925 684.925 -4.595 ;
        RECT 683.235 -4.925 683.565 -4.595 ;
        RECT 681.875 -4.925 682.205 -4.595 ;
        RECT 680.515 -4.925 680.845 -4.595 ;
        RECT 679.155 -4.925 679.485 -4.595 ;
        RECT 678.125 -4.92 954.88 -4.6 ;
        RECT 953.875 -4.925 954.205 -4.595 ;
        RECT 952.515 -4.925 952.845 -4.595 ;
        RECT 951.155 -4.925 951.485 -4.595 ;
        RECT 949.795 -4.925 950.125 -4.595 ;
        RECT 948.435 -4.925 948.765 -4.595 ;
        RECT 947.075 -4.925 947.405 -4.595 ;
        RECT 945.715 -4.925 946.045 -4.595 ;
        RECT 944.355 -4.925 944.685 -4.595 ;
        RECT 942.995 -4.925 943.325 -4.595 ;
        RECT 941.635 -4.925 941.965 -4.595 ;
        RECT 940.275 -4.925 940.605 -4.595 ;
        RECT 938.915 -4.925 939.245 -4.595 ;
        RECT 937.555 -4.925 937.885 -4.595 ;
        RECT 936.195 -4.925 936.525 -4.595 ;
        RECT 934.835 -4.925 935.165 -4.595 ;
        RECT 933.475 -4.925 933.805 -4.595 ;
        RECT 932.115 -4.925 932.445 -4.595 ;
        RECT 930.755 -4.925 931.085 -4.595 ;
        RECT 929.395 -4.925 929.725 -4.595 ;
        RECT 928.035 -4.925 928.365 -4.595 ;
        RECT 926.675 -4.925 927.005 -4.595 ;
        RECT 925.315 -4.925 925.645 -4.595 ;
        RECT 923.955 -4.925 924.285 -4.595 ;
        RECT 922.595 -4.925 922.925 -4.595 ;
        RECT 921.235 -4.925 921.565 -4.595 ;
        RECT 919.875 -4.925 920.205 -4.595 ;
        RECT 918.515 -4.925 918.845 -4.595 ;
        RECT 917.155 -4.925 917.485 -4.595 ;
        RECT 915.795 -4.925 916.125 -4.595 ;
        RECT 914.435 -4.925 914.765 -4.595 ;
        RECT 913.075 -4.925 913.405 -4.595 ;
        RECT 911.715 -4.925 912.045 -4.595 ;
        RECT 910.355 -4.925 910.685 -4.595 ;
        RECT 908.995 -4.925 909.325 -4.595 ;
        RECT 907.635 -4.925 907.965 -4.595 ;
        RECT 906.275 -4.925 906.605 -4.595 ;
        RECT 904.915 -4.925 905.245 -4.595 ;
        RECT 903.555 -4.925 903.885 -4.595 ;
        RECT 902.195 -4.925 902.525 -4.595 ;
        RECT 900.835 -4.925 901.165 -4.595 ;
        RECT 899.475 -4.925 899.805 -4.595 ;
        RECT 898.115 -4.925 898.445 -4.595 ;
        RECT 896.755 -4.925 897.085 -4.595 ;
        RECT 895.395 -4.925 895.725 -4.595 ;
        RECT 894.035 -4.925 894.365 -4.595 ;
        RECT 892.675 -4.925 893.005 -4.595 ;
        RECT 891.315 -4.925 891.645 -4.595 ;
        RECT 889.955 -4.925 890.285 -4.595 ;
        RECT 888.595 -4.925 888.925 -4.595 ;
        RECT 887.235 -4.925 887.565 -4.595 ;
        RECT 885.875 -4.925 886.205 -4.595 ;
        RECT 884.515 -4.925 884.845 -4.595 ;
        RECT 883.155 -4.925 883.485 -4.595 ;
        RECT 881.795 -4.925 882.125 -4.595 ;
        RECT 880.435 -4.925 880.765 -4.595 ;
        RECT 879.075 -4.925 879.405 -4.595 ;
        RECT 877.715 -4.925 878.045 -4.595 ;
        RECT 876.355 -4.925 876.685 -4.595 ;
        RECT 874.995 -4.925 875.325 -4.595 ;
        RECT 873.635 -4.925 873.965 -4.595 ;
        RECT 872.275 -4.925 872.605 -4.595 ;
        RECT 870.915 -4.925 871.245 -4.595 ;
        RECT 869.555 -4.925 869.885 -4.595 ;
        RECT 868.195 -4.925 868.525 -4.595 ;
        RECT 866.835 -4.925 867.165 -4.595 ;
        RECT 865.475 -4.925 865.805 -4.595 ;
        RECT 864.115 -4.925 864.445 -4.595 ;
        RECT 862.755 -4.925 863.085 -4.595 ;
        RECT 861.395 -4.925 861.725 -4.595 ;
        RECT 860.035 -4.925 860.365 -4.595 ;
        RECT 858.675 -4.925 859.005 -4.595 ;
        RECT 857.315 -4.925 857.645 -4.595 ;
        RECT 855.955 -4.925 856.285 -4.595 ;
        RECT 854.595 -4.925 854.925 -4.595 ;
        RECT 853.235 -4.925 853.565 -4.595 ;
        RECT 851.875 -4.925 852.205 -4.595 ;
        RECT 850.515 -4.925 850.845 -4.595 ;
        RECT 849.155 -4.925 849.485 -4.595 ;
        RECT 847.795 -4.925 848.125 -4.595 ;
        RECT 846.435 -4.925 846.765 -4.595 ;
        RECT 845.075 -4.925 845.405 -4.595 ;
        RECT 843.715 -4.925 844.045 -4.595 ;
        RECT 842.355 -4.925 842.685 -4.595 ;
        RECT 840.995 -4.925 841.325 -4.595 ;
        RECT 839.635 -4.925 839.965 -4.595 ;
        RECT 838.275 -4.925 838.605 -4.595 ;
        RECT 836.915 -4.925 837.245 -4.595 ;
        RECT 835.555 -4.925 835.885 -4.595 ;
        RECT 834.195 -4.925 834.525 -4.595 ;
        RECT 832.835 -4.925 833.165 -4.595 ;
        RECT 831.475 -4.925 831.805 -4.595 ;
        RECT 830.115 -4.925 830.445 -4.595 ;
        RECT 828.755 -4.925 829.085 -4.595 ;
        RECT 827.395 -4.925 827.725 -4.595 ;
        RECT 826.035 -4.925 826.365 -4.595 ;
        RECT 824.675 -4.925 825.005 -4.595 ;
        RECT 823.315 -4.925 823.645 -4.595 ;
        RECT 821.955 -4.925 822.285 -4.595 ;
        RECT 820.595 -4.925 820.925 -4.595 ;
        RECT 819.235 -4.925 819.565 -4.595 ;
        RECT 817.875 -4.925 818.205 -4.595 ;
        RECT 816.515 -4.925 816.845 -4.595 ;
        RECT 815.155 -4.925 815.485 -4.595 ;
        RECT 813.795 -4.925 814.125 -4.595 ;
        RECT 812.435 -4.925 812.765 -4.595 ;
        RECT 811.075 -4.925 811.405 -4.595 ;
        RECT 809.715 -4.925 810.045 -4.595 ;
        RECT 808.355 -4.925 808.685 -4.595 ;
        RECT 806.995 -4.925 807.325 -4.595 ;
        RECT 805.635 -4.925 805.965 -4.595 ;
        RECT 804.275 -4.925 804.605 -4.595 ;
        RECT 802.915 -4.925 803.245 -4.595 ;
        RECT 801.555 -4.925 801.885 -4.595 ;
        RECT 800.195 -4.925 800.525 -4.595 ;
        RECT 798.835 -4.925 799.165 -4.595 ;
        RECT 797.475 -4.925 797.805 -4.595 ;
        RECT 796.115 -4.925 796.445 -4.595 ;
        RECT 794.755 -4.925 795.085 -4.595 ;
        RECT 793.395 -4.925 793.725 -4.595 ;
        RECT 792.035 -4.925 792.365 -4.595 ;
        RECT 790.675 -4.925 791.005 -4.595 ;
        RECT 789.315 -4.925 789.645 -4.595 ;
        RECT 787.955 -4.925 788.285 -4.595 ;
        RECT 786.595 -4.925 786.925 -4.595 ;
        RECT 785.235 -4.925 785.565 -4.595 ;
        RECT 783.875 -4.925 784.205 -4.595 ;
        RECT 782.515 -4.925 782.845 -4.595 ;
        RECT 781.155 -4.925 781.485 -4.595 ;
        RECT 779.795 -4.925 780.125 -4.595 ;
        RECT 778.435 -4.925 778.765 -4.595 ;
        RECT 777.075 -4.925 777.405 -4.595 ;
        RECT 775.715 -4.925 776.045 -4.595 ;
        RECT 774.355 -4.925 774.685 -4.595 ;
        RECT 772.995 -4.925 773.325 -4.595 ;
        RECT 771.635 -4.925 771.965 -4.595 ;
        RECT 770.275 -4.925 770.605 -4.595 ;
        RECT 768.915 -4.925 769.245 -4.595 ;
        RECT 767.555 -4.925 767.885 -4.595 ;
        RECT 766.195 -4.925 766.525 -4.595 ;
        RECT 764.835 -4.925 765.165 -4.595 ;
        RECT 763.475 -4.925 763.805 -4.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 -6.285 134.125 -5.955 ;
        RECT 132.435 -6.285 132.765 -5.955 ;
        RECT 131.075 -6.285 131.405 -5.955 ;
        RECT 129.715 -6.285 130.045 -5.955 ;
        RECT 128.355 -6.285 128.685 -5.955 ;
        RECT 126.995 -6.285 127.325 -5.955 ;
        RECT 125.635 -6.285 125.965 -5.955 ;
        RECT 124.275 -6.285 124.605 -5.955 ;
        RECT 122.915 -6.285 123.245 -5.955 ;
        RECT 121.555 -6.285 121.885 -5.955 ;
        RECT 120.195 -6.285 120.525 -5.955 ;
        RECT 118.835 -6.285 119.165 -5.955 ;
        RECT 117.475 -6.285 117.805 -5.955 ;
        RECT 116.115 -6.285 116.445 -5.955 ;
        RECT 114.755 -6.285 115.085 -5.955 ;
        RECT 113.395 -6.285 113.725 -5.955 ;
        RECT 112.035 -6.285 112.365 -5.955 ;
        RECT 110.675 -6.285 111.005 -5.955 ;
        RECT 109.315 -6.285 109.645 -5.955 ;
        RECT 107.955 -6.285 108.285 -5.955 ;
        RECT 106.595 -6.285 106.925 -5.955 ;
        RECT 105.235 -6.285 105.565 -5.955 ;
        RECT 103.875 -6.285 104.205 -5.955 ;
        RECT 102.515 -6.285 102.845 -5.955 ;
        RECT 101.155 -6.285 101.485 -5.955 ;
        RECT 99.795 -6.285 100.125 -5.955 ;
        RECT 98.435 -6.285 98.765 -5.955 ;
        RECT 97.075 -6.285 97.405 -5.955 ;
        RECT 95.715 -6.285 96.045 -5.955 ;
        RECT 94.355 -6.285 94.685 -5.955 ;
        RECT 92.995 -6.285 93.325 -5.955 ;
        RECT 91.635 -6.285 91.965 -5.955 ;
        RECT 90.275 -6.285 90.605 -5.955 ;
        RECT 88.915 -6.285 89.245 -5.955 ;
        RECT 87.555 -6.285 87.885 -5.955 ;
        RECT 86.195 -6.285 86.525 -5.955 ;
        RECT 84.835 -6.285 85.165 -5.955 ;
        RECT 83.475 -6.285 83.805 -5.955 ;
        RECT 82.115 -6.285 82.445 -5.955 ;
        RECT 80.755 -6.285 81.085 -5.955 ;
        RECT 79.395 -6.285 79.725 -5.955 ;
        RECT 78.035 -6.285 78.365 -5.955 ;
        RECT 76.675 -6.285 77.005 -5.955 ;
        RECT 75.315 -6.285 75.645 -5.955 ;
        RECT 73.955 -6.285 74.285 -5.955 ;
        RECT 72.595 -6.285 72.925 -5.955 ;
        RECT 71.235 -6.285 71.565 -5.955 ;
        RECT 69.875 -6.285 70.205 -5.955 ;
        RECT 68.515 -6.285 68.845 -5.955 ;
        RECT 67.155 -6.285 67.485 -5.955 ;
        RECT 65.795 -6.285 66.125 -5.955 ;
        RECT 64.435 -6.285 64.765 -5.955 ;
        RECT 63.075 -6.285 63.405 -5.955 ;
        RECT 61.715 -6.285 62.045 -5.955 ;
        RECT 60.355 -6.285 60.685 -5.955 ;
        RECT 58.995 -6.285 59.325 -5.955 ;
        RECT 57.635 -6.285 57.965 -5.955 ;
        RECT 56.275 -6.285 56.605 -5.955 ;
        RECT 54.915 -6.285 55.245 -5.955 ;
        RECT 53.555 -6.285 53.885 -5.955 ;
        RECT 52.195 -6.285 52.525 -5.955 ;
        RECT 50.835 -6.285 51.165 -5.955 ;
        RECT 49.475 -6.285 49.805 -5.955 ;
        RECT 48.115 -6.285 48.445 -5.955 ;
        RECT 46.755 -6.285 47.085 -5.955 ;
        RECT 45.395 -6.285 45.725 -5.955 ;
        RECT 44.035 -6.285 44.365 -5.955 ;
        RECT 42.675 -6.285 43.005 -5.955 ;
        RECT 41.315 -6.285 41.645 -5.955 ;
        RECT 39.955 -6.285 40.285 -5.955 ;
        RECT 38.595 -6.285 38.925 -5.955 ;
        RECT 37.235 -6.285 37.565 -5.955 ;
        RECT 35.875 -6.285 36.205 -5.955 ;
        RECT 34.515 -6.285 34.845 -5.955 ;
        RECT 33.155 -6.285 33.485 -5.955 ;
        RECT 31.795 -6.285 32.125 -5.955 ;
        RECT 30.435 -6.285 30.765 -5.955 ;
        RECT 29.075 -6.285 29.405 -5.955 ;
        RECT 27.715 -6.285 28.045 -5.955 ;
        RECT 26.355 -6.285 26.685 -5.955 ;
        RECT 24.995 -6.285 25.325 -5.955 ;
        RECT 23.635 -6.285 23.965 -5.955 ;
        RECT 22.275 -6.285 22.605 -5.955 ;
        RECT 20.915 -6.285 21.245 -5.955 ;
        RECT 19.555 -6.285 19.885 -5.955 ;
        RECT 18.195 -6.285 18.525 -5.955 ;
        RECT 16.835 -6.285 17.165 -5.955 ;
        RECT 15.475 -6.285 15.805 -5.955 ;
        RECT 14.115 -6.285 14.445 -5.955 ;
        RECT 12.755 -6.285 13.085 -5.955 ;
        RECT 11.395 -6.285 11.725 -5.955 ;
        RECT 10.035 -6.285 10.365 -5.955 ;
        RECT 8.675 -6.285 9.005 -5.955 ;
        RECT 7.315 -6.285 7.645 -5.955 ;
        RECT 5.955 -6.285 6.285 -5.955 ;
        RECT 4.595 -6.285 4.925 -5.955 ;
        RECT 3.235 -6.285 3.565 -5.955 ;
        RECT 1.875 -6.285 2.205 -5.955 ;
        RECT 0.515 -6.285 0.845 -5.955 ;
        RECT -0.845 -6.285 -0.515 -5.955 ;
        RECT 677.795 -6.285 678.125 -5.955 ;
        RECT -1.52 -6.28 678.125 -5.96 ;
        RECT 676.435 -6.285 676.765 -5.955 ;
        RECT 675.075 -6.285 675.405 -5.955 ;
        RECT 673.715 -6.285 674.045 -5.955 ;
        RECT 672.355 -6.285 672.685 -5.955 ;
        RECT 670.995 -6.285 671.325 -5.955 ;
        RECT 669.635 -6.285 669.965 -5.955 ;
        RECT 668.275 -6.285 668.605 -5.955 ;
        RECT 666.915 -6.285 667.245 -5.955 ;
        RECT 665.555 -6.285 665.885 -5.955 ;
        RECT 664.195 -6.285 664.525 -5.955 ;
        RECT 662.835 -6.285 663.165 -5.955 ;
        RECT 661.475 -6.285 661.805 -5.955 ;
        RECT 660.115 -6.285 660.445 -5.955 ;
        RECT 658.755 -6.285 659.085 -5.955 ;
        RECT 657.395 -6.285 657.725 -5.955 ;
        RECT 656.035 -6.285 656.365 -5.955 ;
        RECT 654.675 -6.285 655.005 -5.955 ;
        RECT 653.315 -6.285 653.645 -5.955 ;
        RECT 651.955 -6.285 652.285 -5.955 ;
        RECT 650.595 -6.285 650.925 -5.955 ;
        RECT 649.235 -6.285 649.565 -5.955 ;
        RECT 647.875 -6.285 648.205 -5.955 ;
        RECT 646.515 -6.285 646.845 -5.955 ;
        RECT 645.155 -6.285 645.485 -5.955 ;
        RECT 643.795 -6.285 644.125 -5.955 ;
        RECT 642.435 -6.285 642.765 -5.955 ;
        RECT 641.075 -6.285 641.405 -5.955 ;
        RECT 639.715 -6.285 640.045 -5.955 ;
        RECT 638.355 -6.285 638.685 -5.955 ;
        RECT 636.995 -6.285 637.325 -5.955 ;
        RECT 635.635 -6.285 635.965 -5.955 ;
        RECT 634.275 -6.285 634.605 -5.955 ;
        RECT 632.915 -6.285 633.245 -5.955 ;
        RECT 631.555 -6.285 631.885 -5.955 ;
        RECT 630.195 -6.285 630.525 -5.955 ;
        RECT 628.835 -6.285 629.165 -5.955 ;
        RECT 627.475 -6.285 627.805 -5.955 ;
        RECT 626.115 -6.285 626.445 -5.955 ;
        RECT 624.755 -6.285 625.085 -5.955 ;
        RECT 623.395 -6.285 623.725 -5.955 ;
        RECT 622.035 -6.285 622.365 -5.955 ;
        RECT 620.675 -6.285 621.005 -5.955 ;
        RECT 619.315 -6.285 619.645 -5.955 ;
        RECT 617.955 -6.285 618.285 -5.955 ;
        RECT 616.595 -6.285 616.925 -5.955 ;
        RECT 615.235 -6.285 615.565 -5.955 ;
        RECT 613.875 -6.285 614.205 -5.955 ;
        RECT 612.515 -6.285 612.845 -5.955 ;
        RECT 611.155 -6.285 611.485 -5.955 ;
        RECT 609.795 -6.285 610.125 -5.955 ;
        RECT 608.435 -6.285 608.765 -5.955 ;
        RECT 607.075 -6.285 607.405 -5.955 ;
        RECT 605.715 -6.285 606.045 -5.955 ;
        RECT 604.355 -6.285 604.685 -5.955 ;
        RECT 602.995 -6.285 603.325 -5.955 ;
        RECT 601.635 -6.285 601.965 -5.955 ;
        RECT 600.275 -6.285 600.605 -5.955 ;
        RECT 598.915 -6.285 599.245 -5.955 ;
        RECT 597.555 -6.285 597.885 -5.955 ;
        RECT 596.195 -6.285 596.525 -5.955 ;
        RECT 594.835 -6.285 595.165 -5.955 ;
        RECT 593.475 -6.285 593.805 -5.955 ;
        RECT 592.115 -6.285 592.445 -5.955 ;
        RECT 590.755 -6.285 591.085 -5.955 ;
        RECT 589.395 -6.285 589.725 -5.955 ;
        RECT 588.035 -6.285 588.365 -5.955 ;
        RECT 586.675 -6.285 587.005 -5.955 ;
        RECT 585.315 -6.285 585.645 -5.955 ;
        RECT 583.955 -6.285 584.285 -5.955 ;
        RECT 582.595 -6.285 582.925 -5.955 ;
        RECT 581.235 -6.285 581.565 -5.955 ;
        RECT 579.875 -6.285 580.205 -5.955 ;
        RECT 578.515 -6.285 578.845 -5.955 ;
        RECT 577.155 -6.285 577.485 -5.955 ;
        RECT 575.795 -6.285 576.125 -5.955 ;
        RECT 574.435 -6.285 574.765 -5.955 ;
        RECT 573.075 -6.285 573.405 -5.955 ;
        RECT 571.715 -6.285 572.045 -5.955 ;
        RECT 570.355 -6.285 570.685 -5.955 ;
        RECT 568.995 -6.285 569.325 -5.955 ;
        RECT 567.635 -6.285 567.965 -5.955 ;
        RECT 566.275 -6.285 566.605 -5.955 ;
        RECT 564.915 -6.285 565.245 -5.955 ;
        RECT 563.555 -6.285 563.885 -5.955 ;
        RECT 562.195 -6.285 562.525 -5.955 ;
        RECT 560.835 -6.285 561.165 -5.955 ;
        RECT 559.475 -6.285 559.805 -5.955 ;
        RECT 558.115 -6.285 558.445 -5.955 ;
        RECT 556.755 -6.285 557.085 -5.955 ;
        RECT 555.395 -6.285 555.725 -5.955 ;
        RECT 554.035 -6.285 554.365 -5.955 ;
        RECT 552.675 -6.285 553.005 -5.955 ;
        RECT 551.315 -6.285 551.645 -5.955 ;
        RECT 549.955 -6.285 550.285 -5.955 ;
        RECT 548.595 -6.285 548.925 -5.955 ;
        RECT 547.235 -6.285 547.565 -5.955 ;
        RECT 545.875 -6.285 546.205 -5.955 ;
        RECT 544.515 -6.285 544.845 -5.955 ;
        RECT 543.155 -6.285 543.485 -5.955 ;
        RECT 541.795 -6.285 542.125 -5.955 ;
        RECT 540.435 -6.285 540.765 -5.955 ;
        RECT 539.075 -6.285 539.405 -5.955 ;
        RECT 537.715 -6.285 538.045 -5.955 ;
        RECT 536.355 -6.285 536.685 -5.955 ;
        RECT 534.995 -6.285 535.325 -5.955 ;
        RECT 533.635 -6.285 533.965 -5.955 ;
        RECT 532.275 -6.285 532.605 -5.955 ;
        RECT 530.915 -6.285 531.245 -5.955 ;
        RECT 529.555 -6.285 529.885 -5.955 ;
        RECT 528.195 -6.285 528.525 -5.955 ;
        RECT 526.835 -6.285 527.165 -5.955 ;
        RECT 525.475 -6.285 525.805 -5.955 ;
        RECT 524.115 -6.285 524.445 -5.955 ;
        RECT 522.755 -6.285 523.085 -5.955 ;
        RECT 521.395 -6.285 521.725 -5.955 ;
        RECT 520.035 -6.285 520.365 -5.955 ;
        RECT 518.675 -6.285 519.005 -5.955 ;
        RECT 517.315 -6.285 517.645 -5.955 ;
        RECT 515.955 -6.285 516.285 -5.955 ;
        RECT 514.595 -6.285 514.925 -5.955 ;
        RECT 513.235 -6.285 513.565 -5.955 ;
        RECT 511.875 -6.285 512.205 -5.955 ;
        RECT 510.515 -6.285 510.845 -5.955 ;
        RECT 509.155 -6.285 509.485 -5.955 ;
        RECT 507.795 -6.285 508.125 -5.955 ;
        RECT 506.435 -6.285 506.765 -5.955 ;
        RECT 505.075 -6.285 505.405 -5.955 ;
        RECT 503.715 -6.285 504.045 -5.955 ;
        RECT 502.355 -6.285 502.685 -5.955 ;
        RECT 500.995 -6.285 501.325 -5.955 ;
        RECT 499.635 -6.285 499.965 -5.955 ;
        RECT 498.275 -6.285 498.605 -5.955 ;
        RECT 496.915 -6.285 497.245 -5.955 ;
        RECT 495.555 -6.285 495.885 -5.955 ;
        RECT 494.195 -6.285 494.525 -5.955 ;
        RECT 492.835 -6.285 493.165 -5.955 ;
        RECT 491.475 -6.285 491.805 -5.955 ;
        RECT 490.115 -6.285 490.445 -5.955 ;
        RECT 488.755 -6.285 489.085 -5.955 ;
        RECT 487.395 -6.285 487.725 -5.955 ;
        RECT 486.035 -6.285 486.365 -5.955 ;
        RECT 484.675 -6.285 485.005 -5.955 ;
        RECT 483.315 -6.285 483.645 -5.955 ;
        RECT 481.955 -6.285 482.285 -5.955 ;
        RECT 480.595 -6.285 480.925 -5.955 ;
        RECT 479.235 -6.285 479.565 -5.955 ;
        RECT 477.875 -6.285 478.205 -5.955 ;
        RECT 476.515 -6.285 476.845 -5.955 ;
        RECT 475.155 -6.285 475.485 -5.955 ;
        RECT 473.795 -6.285 474.125 -5.955 ;
        RECT 472.435 -6.285 472.765 -5.955 ;
        RECT 471.075 -6.285 471.405 -5.955 ;
        RECT 469.715 -6.285 470.045 -5.955 ;
        RECT 468.355 -6.285 468.685 -5.955 ;
        RECT 466.995 -6.285 467.325 -5.955 ;
        RECT 465.635 -6.285 465.965 -5.955 ;
        RECT 464.275 -6.285 464.605 -5.955 ;
        RECT 462.915 -6.285 463.245 -5.955 ;
        RECT 461.555 -6.285 461.885 -5.955 ;
        RECT 460.195 -6.285 460.525 -5.955 ;
        RECT 458.835 -6.285 459.165 -5.955 ;
        RECT 457.475 -6.285 457.805 -5.955 ;
        RECT 456.115 -6.285 456.445 -5.955 ;
        RECT 454.755 -6.285 455.085 -5.955 ;
        RECT 453.395 -6.285 453.725 -5.955 ;
        RECT 452.035 -6.285 452.365 -5.955 ;
        RECT 450.675 -6.285 451.005 -5.955 ;
        RECT 449.315 -6.285 449.645 -5.955 ;
        RECT 447.955 -6.285 448.285 -5.955 ;
        RECT 446.595 -6.285 446.925 -5.955 ;
        RECT 445.235 -6.285 445.565 -5.955 ;
        RECT 443.875 -6.285 444.205 -5.955 ;
        RECT 442.515 -6.285 442.845 -5.955 ;
        RECT 441.155 -6.285 441.485 -5.955 ;
        RECT 439.795 -6.285 440.125 -5.955 ;
        RECT 438.435 -6.285 438.765 -5.955 ;
        RECT 437.075 -6.285 437.405 -5.955 ;
        RECT 435.715 -6.285 436.045 -5.955 ;
        RECT 434.355 -6.285 434.685 -5.955 ;
        RECT 432.995 -6.285 433.325 -5.955 ;
        RECT 431.635 -6.285 431.965 -5.955 ;
        RECT 430.275 -6.285 430.605 -5.955 ;
        RECT 428.915 -6.285 429.245 -5.955 ;
        RECT 427.555 -6.285 427.885 -5.955 ;
        RECT 426.195 -6.285 426.525 -5.955 ;
        RECT 424.835 -6.285 425.165 -5.955 ;
        RECT 423.475 -6.285 423.805 -5.955 ;
        RECT 422.115 -6.285 422.445 -5.955 ;
        RECT 420.755 -6.285 421.085 -5.955 ;
        RECT 419.395 -6.285 419.725 -5.955 ;
        RECT 418.035 -6.285 418.365 -5.955 ;
        RECT 416.675 -6.285 417.005 -5.955 ;
        RECT 415.315 -6.285 415.645 -5.955 ;
        RECT 413.955 -6.285 414.285 -5.955 ;
        RECT 412.595 -6.285 412.925 -5.955 ;
        RECT 411.235 -6.285 411.565 -5.955 ;
        RECT 409.875 -6.285 410.205 -5.955 ;
        RECT 408.515 -6.285 408.845 -5.955 ;
        RECT 407.155 -6.285 407.485 -5.955 ;
        RECT 405.795 -6.285 406.125 -5.955 ;
        RECT 404.435 -6.285 404.765 -5.955 ;
        RECT 403.075 -6.285 403.405 -5.955 ;
        RECT 401.715 -6.285 402.045 -5.955 ;
        RECT 400.355 -6.285 400.685 -5.955 ;
        RECT 398.995 -6.285 399.325 -5.955 ;
        RECT 397.635 -6.285 397.965 -5.955 ;
        RECT 396.275 -6.285 396.605 -5.955 ;
        RECT 394.915 -6.285 395.245 -5.955 ;
        RECT 393.555 -6.285 393.885 -5.955 ;
        RECT 392.195 -6.285 392.525 -5.955 ;
        RECT 390.835 -6.285 391.165 -5.955 ;
        RECT 389.475 -6.285 389.805 -5.955 ;
        RECT 388.115 -6.285 388.445 -5.955 ;
        RECT 386.755 -6.285 387.085 -5.955 ;
        RECT 385.395 -6.285 385.725 -5.955 ;
        RECT 384.035 -6.285 384.365 -5.955 ;
        RECT 382.675 -6.285 383.005 -5.955 ;
        RECT 381.315 -6.285 381.645 -5.955 ;
        RECT 379.955 -6.285 380.285 -5.955 ;
        RECT 378.595 -6.285 378.925 -5.955 ;
        RECT 377.235 -6.285 377.565 -5.955 ;
        RECT 375.875 -6.285 376.205 -5.955 ;
        RECT 374.515 -6.285 374.845 -5.955 ;
        RECT 373.155 -6.285 373.485 -5.955 ;
        RECT 371.795 -6.285 372.125 -5.955 ;
        RECT 370.435 -6.285 370.765 -5.955 ;
        RECT 369.075 -6.285 369.405 -5.955 ;
        RECT 367.715 -6.285 368.045 -5.955 ;
        RECT 366.355 -6.285 366.685 -5.955 ;
        RECT 364.995 -6.285 365.325 -5.955 ;
        RECT 363.635 -6.285 363.965 -5.955 ;
        RECT 362.275 -6.285 362.605 -5.955 ;
        RECT 360.915 -6.285 361.245 -5.955 ;
        RECT 359.555 -6.285 359.885 -5.955 ;
        RECT 358.195 -6.285 358.525 -5.955 ;
        RECT 356.835 -6.285 357.165 -5.955 ;
        RECT 355.475 -6.285 355.805 -5.955 ;
        RECT 354.115 -6.285 354.445 -5.955 ;
        RECT 352.755 -6.285 353.085 -5.955 ;
        RECT 351.395 -6.285 351.725 -5.955 ;
        RECT 350.035 -6.285 350.365 -5.955 ;
        RECT 348.675 -6.285 349.005 -5.955 ;
        RECT 347.315 -6.285 347.645 -5.955 ;
        RECT 345.955 -6.285 346.285 -5.955 ;
        RECT 344.595 -6.285 344.925 -5.955 ;
        RECT 343.235 -6.285 343.565 -5.955 ;
        RECT 341.875 -6.285 342.205 -5.955 ;
        RECT 340.515 -6.285 340.845 -5.955 ;
        RECT 339.155 -6.285 339.485 -5.955 ;
        RECT 337.795 -6.285 338.125 -5.955 ;
        RECT 336.435 -6.285 336.765 -5.955 ;
        RECT 335.075 -6.285 335.405 -5.955 ;
        RECT 333.715 -6.285 334.045 -5.955 ;
        RECT 332.355 -6.285 332.685 -5.955 ;
        RECT 330.995 -6.285 331.325 -5.955 ;
        RECT 329.635 -6.285 329.965 -5.955 ;
        RECT 328.275 -6.285 328.605 -5.955 ;
        RECT 326.915 -6.285 327.245 -5.955 ;
        RECT 325.555 -6.285 325.885 -5.955 ;
        RECT 324.195 -6.285 324.525 -5.955 ;
        RECT 322.835 -6.285 323.165 -5.955 ;
        RECT 321.475 -6.285 321.805 -5.955 ;
        RECT 320.115 -6.285 320.445 -5.955 ;
        RECT 318.755 -6.285 319.085 -5.955 ;
        RECT 317.395 -6.285 317.725 -5.955 ;
        RECT 316.035 -6.285 316.365 -5.955 ;
        RECT 314.675 -6.285 315.005 -5.955 ;
        RECT 313.315 -6.285 313.645 -5.955 ;
        RECT 311.955 -6.285 312.285 -5.955 ;
        RECT 310.595 -6.285 310.925 -5.955 ;
        RECT 309.235 -6.285 309.565 -5.955 ;
        RECT 307.875 -6.285 308.205 -5.955 ;
        RECT 306.515 -6.285 306.845 -5.955 ;
        RECT 305.155 -6.285 305.485 -5.955 ;
        RECT 303.795 -6.285 304.125 -5.955 ;
        RECT 302.435 -6.285 302.765 -5.955 ;
        RECT 301.075 -6.285 301.405 -5.955 ;
        RECT 299.715 -6.285 300.045 -5.955 ;
        RECT 298.355 -6.285 298.685 -5.955 ;
        RECT 296.995 -6.285 297.325 -5.955 ;
        RECT 295.635 -6.285 295.965 -5.955 ;
        RECT 294.275 -6.285 294.605 -5.955 ;
        RECT 292.915 -6.285 293.245 -5.955 ;
        RECT 291.555 -6.285 291.885 -5.955 ;
        RECT 290.195 -6.285 290.525 -5.955 ;
        RECT 288.835 -6.285 289.165 -5.955 ;
        RECT 287.475 -6.285 287.805 -5.955 ;
        RECT 286.115 -6.285 286.445 -5.955 ;
        RECT 284.755 -6.285 285.085 -5.955 ;
        RECT 283.395 -6.285 283.725 -5.955 ;
        RECT 282.035 -6.285 282.365 -5.955 ;
        RECT 280.675 -6.285 281.005 -5.955 ;
        RECT 279.315 -6.285 279.645 -5.955 ;
        RECT 277.955 -6.285 278.285 -5.955 ;
        RECT 276.595 -6.285 276.925 -5.955 ;
        RECT 275.235 -6.285 275.565 -5.955 ;
        RECT 273.875 -6.285 274.205 -5.955 ;
        RECT 272.515 -6.285 272.845 -5.955 ;
        RECT 271.155 -6.285 271.485 -5.955 ;
        RECT 269.795 -6.285 270.125 -5.955 ;
        RECT 268.435 -6.285 268.765 -5.955 ;
        RECT 267.075 -6.285 267.405 -5.955 ;
        RECT 265.715 -6.285 266.045 -5.955 ;
        RECT 264.355 -6.285 264.685 -5.955 ;
        RECT 262.995 -6.285 263.325 -5.955 ;
        RECT 261.635 -6.285 261.965 -5.955 ;
        RECT 260.275 -6.285 260.605 -5.955 ;
        RECT 258.915 -6.285 259.245 -5.955 ;
        RECT 257.555 -6.285 257.885 -5.955 ;
        RECT 256.195 -6.285 256.525 -5.955 ;
        RECT 254.835 -6.285 255.165 -5.955 ;
        RECT 253.475 -6.285 253.805 -5.955 ;
        RECT 252.115 -6.285 252.445 -5.955 ;
        RECT 250.755 -6.285 251.085 -5.955 ;
        RECT 249.395 -6.285 249.725 -5.955 ;
        RECT 248.035 -6.285 248.365 -5.955 ;
        RECT 246.675 -6.285 247.005 -5.955 ;
        RECT 245.315 -6.285 245.645 -5.955 ;
        RECT 243.955 -6.285 244.285 -5.955 ;
        RECT 242.595 -6.285 242.925 -5.955 ;
        RECT 241.235 -6.285 241.565 -5.955 ;
        RECT 239.875 -6.285 240.205 -5.955 ;
        RECT 238.515 -6.285 238.845 -5.955 ;
        RECT 237.155 -6.285 237.485 -5.955 ;
        RECT 235.795 -6.285 236.125 -5.955 ;
        RECT 234.435 -6.285 234.765 -5.955 ;
        RECT 233.075 -6.285 233.405 -5.955 ;
        RECT 231.715 -6.285 232.045 -5.955 ;
        RECT 230.355 -6.285 230.685 -5.955 ;
        RECT 228.995 -6.285 229.325 -5.955 ;
        RECT 227.635 -6.285 227.965 -5.955 ;
        RECT 226.275 -6.285 226.605 -5.955 ;
        RECT 224.915 -6.285 225.245 -5.955 ;
        RECT 223.555 -6.285 223.885 -5.955 ;
        RECT 222.195 -6.285 222.525 -5.955 ;
        RECT 220.835 -6.285 221.165 -5.955 ;
        RECT 219.475 -6.285 219.805 -5.955 ;
        RECT 218.115 -6.285 218.445 -5.955 ;
        RECT 216.755 -6.285 217.085 -5.955 ;
        RECT 215.395 -6.285 215.725 -5.955 ;
        RECT 214.035 -6.285 214.365 -5.955 ;
        RECT 212.675 -6.285 213.005 -5.955 ;
        RECT 211.315 -6.285 211.645 -5.955 ;
        RECT 209.955 -6.285 210.285 -5.955 ;
        RECT 208.595 -6.285 208.925 -5.955 ;
        RECT 207.235 -6.285 207.565 -5.955 ;
        RECT 205.875 -6.285 206.205 -5.955 ;
        RECT 204.515 -6.285 204.845 -5.955 ;
        RECT 203.155 -6.285 203.485 -5.955 ;
        RECT 201.795 -6.285 202.125 -5.955 ;
        RECT 200.435 -6.285 200.765 -5.955 ;
        RECT 199.075 -6.285 199.405 -5.955 ;
        RECT 197.715 -6.285 198.045 -5.955 ;
        RECT 196.355 -6.285 196.685 -5.955 ;
        RECT 194.995 -6.285 195.325 -5.955 ;
        RECT 193.635 -6.285 193.965 -5.955 ;
        RECT 192.275 -6.285 192.605 -5.955 ;
        RECT 190.915 -6.285 191.245 -5.955 ;
        RECT 189.555 -6.285 189.885 -5.955 ;
        RECT 188.195 -6.285 188.525 -5.955 ;
        RECT 186.835 -6.285 187.165 -5.955 ;
        RECT 185.475 -6.285 185.805 -5.955 ;
        RECT 184.115 -6.285 184.445 -5.955 ;
        RECT 182.755 -6.285 183.085 -5.955 ;
        RECT 181.395 -6.285 181.725 -5.955 ;
        RECT 180.035 -6.285 180.365 -5.955 ;
        RECT 178.675 -6.285 179.005 -5.955 ;
        RECT 177.315 -6.285 177.645 -5.955 ;
        RECT 175.955 -6.285 176.285 -5.955 ;
        RECT 174.595 -6.285 174.925 -5.955 ;
        RECT 173.235 -6.285 173.565 -5.955 ;
        RECT 171.875 -6.285 172.205 -5.955 ;
        RECT 170.515 -6.285 170.845 -5.955 ;
        RECT 169.155 -6.285 169.485 -5.955 ;
        RECT 167.795 -6.285 168.125 -5.955 ;
        RECT 166.435 -6.285 166.765 -5.955 ;
        RECT 165.075 -6.285 165.405 -5.955 ;
        RECT 163.715 -6.285 164.045 -5.955 ;
        RECT 162.355 -6.285 162.685 -5.955 ;
        RECT 160.995 -6.285 161.325 -5.955 ;
        RECT 159.635 -6.285 159.965 -5.955 ;
        RECT 158.275 -6.285 158.605 -5.955 ;
        RECT 156.915 -6.285 157.245 -5.955 ;
        RECT 155.555 -6.285 155.885 -5.955 ;
        RECT 154.195 -6.285 154.525 -5.955 ;
        RECT 152.835 -6.285 153.165 -5.955 ;
        RECT 151.475 -6.285 151.805 -5.955 ;
        RECT 150.115 -6.285 150.445 -5.955 ;
        RECT 148.755 -6.285 149.085 -5.955 ;
        RECT 147.395 -6.285 147.725 -5.955 ;
        RECT 146.035 -6.285 146.365 -5.955 ;
        RECT 144.675 -6.285 145.005 -5.955 ;
        RECT 143.315 -6.285 143.645 -5.955 ;
        RECT 141.955 -6.285 142.285 -5.955 ;
        RECT 140.595 -6.285 140.925 -5.955 ;
        RECT 139.235 -6.285 139.565 -5.955 ;
        RECT 137.875 -6.285 138.205 -5.955 ;
        RECT 136.515 -6.285 136.845 -5.955 ;
        RECT 135.155 -6.285 135.485 -5.955 ;
        RECT 678.125 -6.28 954.88 -5.96 ;
        RECT 953.875 -6.285 954.205 -5.955 ;
        RECT 952.515 -6.285 952.845 -5.955 ;
        RECT 951.155 -6.285 951.485 -5.955 ;
        RECT 949.795 -6.285 950.125 -5.955 ;
        RECT 948.435 -6.285 948.765 -5.955 ;
        RECT 947.075 -6.285 947.405 -5.955 ;
        RECT 945.715 -6.285 946.045 -5.955 ;
        RECT 944.355 -6.285 944.685 -5.955 ;
        RECT 942.995 -6.285 943.325 -5.955 ;
        RECT 941.635 -6.285 941.965 -5.955 ;
        RECT 940.275 -6.285 940.605 -5.955 ;
        RECT 938.915 -6.285 939.245 -5.955 ;
        RECT 937.555 -6.285 937.885 -5.955 ;
        RECT 936.195 -6.285 936.525 -5.955 ;
        RECT 934.835 -6.285 935.165 -5.955 ;
        RECT 933.475 -6.285 933.805 -5.955 ;
        RECT 932.115 -6.285 932.445 -5.955 ;
        RECT 930.755 -6.285 931.085 -5.955 ;
        RECT 929.395 -6.285 929.725 -5.955 ;
        RECT 928.035 -6.285 928.365 -5.955 ;
        RECT 926.675 -6.285 927.005 -5.955 ;
        RECT 925.315 -6.285 925.645 -5.955 ;
        RECT 923.955 -6.285 924.285 -5.955 ;
        RECT 922.595 -6.285 922.925 -5.955 ;
        RECT 921.235 -6.285 921.565 -5.955 ;
        RECT 919.875 -6.285 920.205 -5.955 ;
        RECT 918.515 -6.285 918.845 -5.955 ;
        RECT 917.155 -6.285 917.485 -5.955 ;
        RECT 915.795 -6.285 916.125 -5.955 ;
        RECT 914.435 -6.285 914.765 -5.955 ;
        RECT 913.075 -6.285 913.405 -5.955 ;
        RECT 911.715 -6.285 912.045 -5.955 ;
        RECT 910.355 -6.285 910.685 -5.955 ;
        RECT 908.995 -6.285 909.325 -5.955 ;
        RECT 907.635 -6.285 907.965 -5.955 ;
        RECT 906.275 -6.285 906.605 -5.955 ;
        RECT 904.915 -6.285 905.245 -5.955 ;
        RECT 903.555 -6.285 903.885 -5.955 ;
        RECT 902.195 -6.285 902.525 -5.955 ;
        RECT 900.835 -6.285 901.165 -5.955 ;
        RECT 899.475 -6.285 899.805 -5.955 ;
        RECT 898.115 -6.285 898.445 -5.955 ;
        RECT 896.755 -6.285 897.085 -5.955 ;
        RECT 895.395 -6.285 895.725 -5.955 ;
        RECT 894.035 -6.285 894.365 -5.955 ;
        RECT 892.675 -6.285 893.005 -5.955 ;
        RECT 891.315 -6.285 891.645 -5.955 ;
        RECT 889.955 -6.285 890.285 -5.955 ;
        RECT 888.595 -6.285 888.925 -5.955 ;
        RECT 887.235 -6.285 887.565 -5.955 ;
        RECT 885.875 -6.285 886.205 -5.955 ;
        RECT 884.515 -6.285 884.845 -5.955 ;
        RECT 883.155 -6.285 883.485 -5.955 ;
        RECT 881.795 -6.285 882.125 -5.955 ;
        RECT 880.435 -6.285 880.765 -5.955 ;
        RECT 879.075 -6.285 879.405 -5.955 ;
        RECT 877.715 -6.285 878.045 -5.955 ;
        RECT 876.355 -6.285 876.685 -5.955 ;
        RECT 874.995 -6.285 875.325 -5.955 ;
        RECT 873.635 -6.285 873.965 -5.955 ;
        RECT 872.275 -6.285 872.605 -5.955 ;
        RECT 870.915 -6.285 871.245 -5.955 ;
        RECT 869.555 -6.285 869.885 -5.955 ;
        RECT 868.195 -6.285 868.525 -5.955 ;
        RECT 866.835 -6.285 867.165 -5.955 ;
        RECT 865.475 -6.285 865.805 -5.955 ;
        RECT 864.115 -6.285 864.445 -5.955 ;
        RECT 862.755 -6.285 863.085 -5.955 ;
        RECT 861.395 -6.285 861.725 -5.955 ;
        RECT 860.035 -6.285 860.365 -5.955 ;
        RECT 858.675 -6.285 859.005 -5.955 ;
        RECT 857.315 -6.285 857.645 -5.955 ;
        RECT 855.955 -6.285 856.285 -5.955 ;
        RECT 854.595 -6.285 854.925 -5.955 ;
        RECT 853.235 -6.285 853.565 -5.955 ;
        RECT 851.875 -6.285 852.205 -5.955 ;
        RECT 850.515 -6.285 850.845 -5.955 ;
        RECT 849.155 -6.285 849.485 -5.955 ;
        RECT 847.795 -6.285 848.125 -5.955 ;
        RECT 846.435 -6.285 846.765 -5.955 ;
        RECT 845.075 -6.285 845.405 -5.955 ;
        RECT 843.715 -6.285 844.045 -5.955 ;
        RECT 842.355 -6.285 842.685 -5.955 ;
        RECT 840.995 -6.285 841.325 -5.955 ;
        RECT 839.635 -6.285 839.965 -5.955 ;
        RECT 838.275 -6.285 838.605 -5.955 ;
        RECT 836.915 -6.285 837.245 -5.955 ;
        RECT 835.555 -6.285 835.885 -5.955 ;
        RECT 834.195 -6.285 834.525 -5.955 ;
        RECT 832.835 -6.285 833.165 -5.955 ;
        RECT 831.475 -6.285 831.805 -5.955 ;
        RECT 830.115 -6.285 830.445 -5.955 ;
        RECT 828.755 -6.285 829.085 -5.955 ;
        RECT 827.395 -6.285 827.725 -5.955 ;
        RECT 826.035 -6.285 826.365 -5.955 ;
        RECT 824.675 -6.285 825.005 -5.955 ;
        RECT 823.315 -6.285 823.645 -5.955 ;
        RECT 821.955 -6.285 822.285 -5.955 ;
        RECT 820.595 -6.285 820.925 -5.955 ;
        RECT 819.235 -6.285 819.565 -5.955 ;
        RECT 817.875 -6.285 818.205 -5.955 ;
        RECT 816.515 -6.285 816.845 -5.955 ;
        RECT 815.155 -6.285 815.485 -5.955 ;
        RECT 813.795 -6.285 814.125 -5.955 ;
        RECT 812.435 -6.285 812.765 -5.955 ;
        RECT 811.075 -6.285 811.405 -5.955 ;
        RECT 809.715 -6.285 810.045 -5.955 ;
        RECT 808.355 -6.285 808.685 -5.955 ;
        RECT 806.995 -6.285 807.325 -5.955 ;
        RECT 805.635 -6.285 805.965 -5.955 ;
        RECT 804.275 -6.285 804.605 -5.955 ;
        RECT 802.915 -6.285 803.245 -5.955 ;
        RECT 801.555 -6.285 801.885 -5.955 ;
        RECT 800.195 -6.285 800.525 -5.955 ;
        RECT 798.835 -6.285 799.165 -5.955 ;
        RECT 797.475 -6.285 797.805 -5.955 ;
        RECT 796.115 -6.285 796.445 -5.955 ;
        RECT 794.755 -6.285 795.085 -5.955 ;
        RECT 793.395 -6.285 793.725 -5.955 ;
        RECT 792.035 -6.285 792.365 -5.955 ;
        RECT 790.675 -6.285 791.005 -5.955 ;
        RECT 789.315 -6.285 789.645 -5.955 ;
        RECT 787.955 -6.285 788.285 -5.955 ;
        RECT 786.595 -6.285 786.925 -5.955 ;
        RECT 785.235 -6.285 785.565 -5.955 ;
        RECT 783.875 -6.285 784.205 -5.955 ;
        RECT 782.515 -6.285 782.845 -5.955 ;
        RECT 781.155 -6.285 781.485 -5.955 ;
        RECT 779.795 -6.285 780.125 -5.955 ;
        RECT 778.435 -6.285 778.765 -5.955 ;
        RECT 777.075 -6.285 777.405 -5.955 ;
        RECT 775.715 -6.285 776.045 -5.955 ;
        RECT 774.355 -6.285 774.685 -5.955 ;
        RECT 772.995 -6.285 773.325 -5.955 ;
        RECT 771.635 -6.285 771.965 -5.955 ;
        RECT 770.275 -6.285 770.605 -5.955 ;
        RECT 768.915 -6.285 769.245 -5.955 ;
        RECT 767.555 -6.285 767.885 -5.955 ;
        RECT 766.195 -6.285 766.525 -5.955 ;
        RECT 764.835 -6.285 765.165 -5.955 ;
        RECT 763.475 -6.285 763.805 -5.955 ;
        RECT 762.115 -6.285 762.445 -5.955 ;
        RECT 760.755 -6.285 761.085 -5.955 ;
        RECT 759.395 -6.285 759.725 -5.955 ;
        RECT 758.035 -6.285 758.365 -5.955 ;
        RECT 756.675 -6.285 757.005 -5.955 ;
        RECT 755.315 -6.285 755.645 -5.955 ;
        RECT 753.955 -6.285 754.285 -5.955 ;
        RECT 752.595 -6.285 752.925 -5.955 ;
        RECT 751.235 -6.285 751.565 -5.955 ;
        RECT 749.875 -6.285 750.205 -5.955 ;
        RECT 748.515 -6.285 748.845 -5.955 ;
        RECT 747.155 -6.285 747.485 -5.955 ;
        RECT 745.795 -6.285 746.125 -5.955 ;
        RECT 744.435 -6.285 744.765 -5.955 ;
        RECT 743.075 -6.285 743.405 -5.955 ;
        RECT 741.715 -6.285 742.045 -5.955 ;
        RECT 740.355 -6.285 740.685 -5.955 ;
        RECT 738.995 -6.285 739.325 -5.955 ;
        RECT 737.635 -6.285 737.965 -5.955 ;
        RECT 736.275 -6.285 736.605 -5.955 ;
        RECT 734.915 -6.285 735.245 -5.955 ;
        RECT 733.555 -6.285 733.885 -5.955 ;
        RECT 732.195 -6.285 732.525 -5.955 ;
        RECT 730.835 -6.285 731.165 -5.955 ;
        RECT 729.475 -6.285 729.805 -5.955 ;
        RECT 728.115 -6.285 728.445 -5.955 ;
        RECT 726.755 -6.285 727.085 -5.955 ;
        RECT 725.395 -6.285 725.725 -5.955 ;
        RECT 724.035 -6.285 724.365 -5.955 ;
        RECT 722.675 -6.285 723.005 -5.955 ;
        RECT 721.315 -6.285 721.645 -5.955 ;
        RECT 719.955 -6.285 720.285 -5.955 ;
        RECT 718.595 -6.285 718.925 -5.955 ;
        RECT 717.235 -6.285 717.565 -5.955 ;
        RECT 715.875 -6.285 716.205 -5.955 ;
        RECT 714.515 -6.285 714.845 -5.955 ;
        RECT 713.155 -6.285 713.485 -5.955 ;
        RECT 711.795 -6.285 712.125 -5.955 ;
        RECT 710.435 -6.285 710.765 -5.955 ;
        RECT 709.075 -6.285 709.405 -5.955 ;
        RECT 707.715 -6.285 708.045 -5.955 ;
        RECT 706.355 -6.285 706.685 -5.955 ;
        RECT 704.995 -6.285 705.325 -5.955 ;
        RECT 703.635 -6.285 703.965 -5.955 ;
        RECT 702.275 -6.285 702.605 -5.955 ;
        RECT 700.915 -6.285 701.245 -5.955 ;
        RECT 699.555 -6.285 699.885 -5.955 ;
        RECT 698.195 -6.285 698.525 -5.955 ;
        RECT 696.835 -6.285 697.165 -5.955 ;
        RECT 695.475 -6.285 695.805 -5.955 ;
        RECT 694.115 -6.285 694.445 -5.955 ;
        RECT 692.755 -6.285 693.085 -5.955 ;
        RECT 691.395 -6.285 691.725 -5.955 ;
        RECT 690.035 -6.285 690.365 -5.955 ;
        RECT 688.675 -6.285 689.005 -5.955 ;
        RECT 687.315 -6.285 687.645 -5.955 ;
        RECT 685.955 -6.285 686.285 -5.955 ;
        RECT 684.595 -6.285 684.925 -5.955 ;
        RECT 683.235 -6.285 683.565 -5.955 ;
        RECT 681.875 -6.285 682.205 -5.955 ;
        RECT 680.515 -6.285 680.845 -5.955 ;
        RECT 679.155 -6.285 679.485 -5.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 -2.205 678.125 -1.875 ;
        RECT -1.52 -2.2 678.125 -1.88 ;
        RECT 676.435 -2.205 676.765 -1.875 ;
        RECT 675.075 -2.205 675.405 -1.875 ;
        RECT 673.715 -2.205 674.045 -1.875 ;
        RECT 672.355 -2.205 672.685 -1.875 ;
        RECT 670.995 -2.205 671.325 -1.875 ;
        RECT 669.635 -2.205 669.965 -1.875 ;
        RECT 668.275 -2.205 668.605 -1.875 ;
        RECT 666.915 -2.205 667.245 -1.875 ;
        RECT 665.555 -2.205 665.885 -1.875 ;
        RECT 664.195 -2.205 664.525 -1.875 ;
        RECT 662.835 -2.205 663.165 -1.875 ;
        RECT 661.475 -2.205 661.805 -1.875 ;
        RECT 660.115 -2.205 660.445 -1.875 ;
        RECT 658.755 -2.205 659.085 -1.875 ;
        RECT 657.395 -2.205 657.725 -1.875 ;
        RECT 656.035 -2.205 656.365 -1.875 ;
        RECT 654.675 -2.205 655.005 -1.875 ;
        RECT 653.315 -2.205 653.645 -1.875 ;
        RECT 651.955 -2.205 652.285 -1.875 ;
        RECT 650.595 -2.205 650.925 -1.875 ;
        RECT 649.235 -2.205 649.565 -1.875 ;
        RECT 647.875 -2.205 648.205 -1.875 ;
        RECT 646.515 -2.205 646.845 -1.875 ;
        RECT 645.155 -2.205 645.485 -1.875 ;
        RECT 643.795 -2.205 644.125 -1.875 ;
        RECT 642.435 -2.205 642.765 -1.875 ;
        RECT 641.075 -2.205 641.405 -1.875 ;
        RECT 639.715 -2.205 640.045 -1.875 ;
        RECT 638.355 -2.205 638.685 -1.875 ;
        RECT 636.995 -2.205 637.325 -1.875 ;
        RECT 635.635 -2.205 635.965 -1.875 ;
        RECT 634.275 -2.205 634.605 -1.875 ;
        RECT 632.915 -2.205 633.245 -1.875 ;
        RECT 631.555 -2.205 631.885 -1.875 ;
        RECT 630.195 -2.205 630.525 -1.875 ;
        RECT 628.835 -2.205 629.165 -1.875 ;
        RECT 627.475 -2.205 627.805 -1.875 ;
        RECT 626.115 -2.205 626.445 -1.875 ;
        RECT 624.755 -2.205 625.085 -1.875 ;
        RECT 623.395 -2.205 623.725 -1.875 ;
        RECT 622.035 -2.205 622.365 -1.875 ;
        RECT 620.675 -2.205 621.005 -1.875 ;
        RECT 619.315 -2.205 619.645 -1.875 ;
        RECT 617.955 -2.205 618.285 -1.875 ;
        RECT 616.595 -2.205 616.925 -1.875 ;
        RECT 615.235 -2.205 615.565 -1.875 ;
        RECT 613.875 -2.205 614.205 -1.875 ;
        RECT 612.515 -2.205 612.845 -1.875 ;
        RECT 611.155 -2.205 611.485 -1.875 ;
        RECT 609.795 -2.205 610.125 -1.875 ;
        RECT 608.435 -2.205 608.765 -1.875 ;
        RECT 607.075 -2.205 607.405 -1.875 ;
        RECT 605.715 -2.205 606.045 -1.875 ;
        RECT 604.355 -2.205 604.685 -1.875 ;
        RECT 602.995 -2.205 603.325 -1.875 ;
        RECT 601.635 -2.205 601.965 -1.875 ;
        RECT 600.275 -2.205 600.605 -1.875 ;
        RECT 598.915 -2.205 599.245 -1.875 ;
        RECT 597.555 -2.205 597.885 -1.875 ;
        RECT 596.195 -2.205 596.525 -1.875 ;
        RECT 594.835 -2.205 595.165 -1.875 ;
        RECT 593.475 -2.205 593.805 -1.875 ;
        RECT 592.115 -2.205 592.445 -1.875 ;
        RECT 590.755 -2.205 591.085 -1.875 ;
        RECT 589.395 -2.205 589.725 -1.875 ;
        RECT 588.035 -2.205 588.365 -1.875 ;
        RECT 586.675 -2.205 587.005 -1.875 ;
        RECT 585.315 -2.205 585.645 -1.875 ;
        RECT 583.955 -2.205 584.285 -1.875 ;
        RECT 582.595 -2.205 582.925 -1.875 ;
        RECT 581.235 -2.205 581.565 -1.875 ;
        RECT 579.875 -2.205 580.205 -1.875 ;
        RECT 578.515 -2.205 578.845 -1.875 ;
        RECT 577.155 -2.205 577.485 -1.875 ;
        RECT 575.795 -2.205 576.125 -1.875 ;
        RECT 574.435 -2.205 574.765 -1.875 ;
        RECT 573.075 -2.205 573.405 -1.875 ;
        RECT 571.715 -2.205 572.045 -1.875 ;
        RECT 570.355 -2.205 570.685 -1.875 ;
        RECT 568.995 -2.205 569.325 -1.875 ;
        RECT 567.635 -2.205 567.965 -1.875 ;
        RECT 566.275 -2.205 566.605 -1.875 ;
        RECT 564.915 -2.205 565.245 -1.875 ;
        RECT 563.555 -2.205 563.885 -1.875 ;
        RECT 562.195 -2.205 562.525 -1.875 ;
        RECT 560.835 -2.205 561.165 -1.875 ;
        RECT 559.475 -2.205 559.805 -1.875 ;
        RECT 558.115 -2.205 558.445 -1.875 ;
        RECT 556.755 -2.205 557.085 -1.875 ;
        RECT 555.395 -2.205 555.725 -1.875 ;
        RECT 554.035 -2.205 554.365 -1.875 ;
        RECT 552.675 -2.205 553.005 -1.875 ;
        RECT 551.315 -2.205 551.645 -1.875 ;
        RECT 549.955 -2.205 550.285 -1.875 ;
        RECT 548.595 -2.205 548.925 -1.875 ;
        RECT 547.235 -2.205 547.565 -1.875 ;
        RECT 545.875 -2.205 546.205 -1.875 ;
        RECT 544.515 -2.205 544.845 -1.875 ;
        RECT 543.155 -2.205 543.485 -1.875 ;
        RECT 541.795 -2.205 542.125 -1.875 ;
        RECT 540.435 -2.205 540.765 -1.875 ;
        RECT 539.075 -2.205 539.405 -1.875 ;
        RECT 537.715 -2.205 538.045 -1.875 ;
        RECT 536.355 -2.205 536.685 -1.875 ;
        RECT 534.995 -2.205 535.325 -1.875 ;
        RECT 533.635 -2.205 533.965 -1.875 ;
        RECT 532.275 -2.205 532.605 -1.875 ;
        RECT 530.915 -2.205 531.245 -1.875 ;
        RECT 529.555 -2.205 529.885 -1.875 ;
        RECT 528.195 -2.205 528.525 -1.875 ;
        RECT 526.835 -2.205 527.165 -1.875 ;
        RECT 525.475 -2.205 525.805 -1.875 ;
        RECT 524.115 -2.205 524.445 -1.875 ;
        RECT 522.755 -2.205 523.085 -1.875 ;
        RECT 521.395 -2.205 521.725 -1.875 ;
        RECT 520.035 -2.205 520.365 -1.875 ;
        RECT 518.675 -2.205 519.005 -1.875 ;
        RECT 517.315 -2.205 517.645 -1.875 ;
        RECT 515.955 -2.205 516.285 -1.875 ;
        RECT 514.595 -2.205 514.925 -1.875 ;
        RECT 513.235 -2.205 513.565 -1.875 ;
        RECT 511.875 -2.205 512.205 -1.875 ;
        RECT 510.515 -2.205 510.845 -1.875 ;
        RECT 509.155 -2.205 509.485 -1.875 ;
        RECT 507.795 -2.205 508.125 -1.875 ;
        RECT 506.435 -2.205 506.765 -1.875 ;
        RECT 505.075 -2.205 505.405 -1.875 ;
        RECT 503.715 -2.205 504.045 -1.875 ;
        RECT 502.355 -2.205 502.685 -1.875 ;
        RECT 500.995 -2.205 501.325 -1.875 ;
        RECT 499.635 -2.205 499.965 -1.875 ;
        RECT 498.275 -2.205 498.605 -1.875 ;
        RECT 496.915 -2.205 497.245 -1.875 ;
        RECT 495.555 -2.205 495.885 -1.875 ;
        RECT 494.195 -2.205 494.525 -1.875 ;
        RECT 492.835 -2.205 493.165 -1.875 ;
        RECT 491.475 -2.205 491.805 -1.875 ;
        RECT 490.115 -2.205 490.445 -1.875 ;
        RECT 488.755 -2.205 489.085 -1.875 ;
        RECT 487.395 -2.205 487.725 -1.875 ;
        RECT 486.035 -2.205 486.365 -1.875 ;
        RECT 484.675 -2.205 485.005 -1.875 ;
        RECT 483.315 -2.205 483.645 -1.875 ;
        RECT 481.955 -2.205 482.285 -1.875 ;
        RECT 480.595 -2.205 480.925 -1.875 ;
        RECT 479.235 -2.205 479.565 -1.875 ;
        RECT 477.875 -2.205 478.205 -1.875 ;
        RECT 476.515 -2.205 476.845 -1.875 ;
        RECT 475.155 -2.205 475.485 -1.875 ;
        RECT 473.795 -2.205 474.125 -1.875 ;
        RECT 472.435 -2.205 472.765 -1.875 ;
        RECT 471.075 -2.205 471.405 -1.875 ;
        RECT 469.715 -2.205 470.045 -1.875 ;
        RECT 468.355 -2.205 468.685 -1.875 ;
        RECT 466.995 -2.205 467.325 -1.875 ;
        RECT 465.635 -2.205 465.965 -1.875 ;
        RECT 464.275 -2.205 464.605 -1.875 ;
        RECT 462.915 -2.205 463.245 -1.875 ;
        RECT 461.555 -2.205 461.885 -1.875 ;
        RECT 460.195 -2.205 460.525 -1.875 ;
        RECT 458.835 -2.205 459.165 -1.875 ;
        RECT 457.475 -2.205 457.805 -1.875 ;
        RECT 456.115 -2.205 456.445 -1.875 ;
        RECT 454.755 -2.205 455.085 -1.875 ;
        RECT 453.395 -2.205 453.725 -1.875 ;
        RECT 452.035 -2.205 452.365 -1.875 ;
        RECT 450.675 -2.205 451.005 -1.875 ;
        RECT 449.315 -2.205 449.645 -1.875 ;
        RECT 447.955 -2.205 448.285 -1.875 ;
        RECT 446.595 -2.205 446.925 -1.875 ;
        RECT 445.235 -2.205 445.565 -1.875 ;
        RECT 443.875 -2.205 444.205 -1.875 ;
        RECT 442.515 -2.205 442.845 -1.875 ;
        RECT 441.155 -2.205 441.485 -1.875 ;
        RECT 439.795 -2.205 440.125 -1.875 ;
        RECT 438.435 -2.205 438.765 -1.875 ;
        RECT 437.075 -2.205 437.405 -1.875 ;
        RECT 435.715 -2.205 436.045 -1.875 ;
        RECT 434.355 -2.205 434.685 -1.875 ;
        RECT 432.995 -2.205 433.325 -1.875 ;
        RECT 431.635 -2.205 431.965 -1.875 ;
        RECT 430.275 -2.205 430.605 -1.875 ;
        RECT 428.915 -2.205 429.245 -1.875 ;
        RECT 427.555 -2.205 427.885 -1.875 ;
        RECT 426.195 -2.205 426.525 -1.875 ;
        RECT 424.835 -2.205 425.165 -1.875 ;
        RECT 423.475 -2.205 423.805 -1.875 ;
        RECT 422.115 -2.205 422.445 -1.875 ;
        RECT 420.755 -2.205 421.085 -1.875 ;
        RECT 419.395 -2.205 419.725 -1.875 ;
        RECT 418.035 -2.205 418.365 -1.875 ;
        RECT 416.675 -2.205 417.005 -1.875 ;
        RECT 415.315 -2.205 415.645 -1.875 ;
        RECT 413.955 -2.205 414.285 -1.875 ;
        RECT 412.595 -2.205 412.925 -1.875 ;
        RECT 411.235 -2.205 411.565 -1.875 ;
        RECT 409.875 -2.205 410.205 -1.875 ;
        RECT 408.515 -2.205 408.845 -1.875 ;
        RECT 407.155 -2.205 407.485 -1.875 ;
        RECT 405.795 -2.205 406.125 -1.875 ;
        RECT 404.435 -2.205 404.765 -1.875 ;
        RECT 403.075 -2.205 403.405 -1.875 ;
        RECT 401.715 -2.205 402.045 -1.875 ;
        RECT 400.355 -2.205 400.685 -1.875 ;
        RECT 398.995 -2.205 399.325 -1.875 ;
        RECT 397.635 -2.205 397.965 -1.875 ;
        RECT 396.275 -2.205 396.605 -1.875 ;
        RECT 394.915 -2.205 395.245 -1.875 ;
        RECT 393.555 -2.205 393.885 -1.875 ;
        RECT 392.195 -2.205 392.525 -1.875 ;
        RECT 390.835 -2.205 391.165 -1.875 ;
        RECT 389.475 -2.205 389.805 -1.875 ;
        RECT 388.115 -2.205 388.445 -1.875 ;
        RECT 386.755 -2.205 387.085 -1.875 ;
        RECT 385.395 -2.205 385.725 -1.875 ;
        RECT 384.035 -2.205 384.365 -1.875 ;
        RECT 382.675 -2.205 383.005 -1.875 ;
        RECT 381.315 -2.205 381.645 -1.875 ;
        RECT 379.955 -2.205 380.285 -1.875 ;
        RECT 378.595 -2.205 378.925 -1.875 ;
        RECT 377.235 -2.205 377.565 -1.875 ;
        RECT 375.875 -2.205 376.205 -1.875 ;
        RECT 374.515 -2.205 374.845 -1.875 ;
        RECT 373.155 -2.205 373.485 -1.875 ;
        RECT 371.795 -2.205 372.125 -1.875 ;
        RECT 370.435 -2.205 370.765 -1.875 ;
        RECT 369.075 -2.205 369.405 -1.875 ;
        RECT 367.715 -2.205 368.045 -1.875 ;
        RECT 366.355 -2.205 366.685 -1.875 ;
        RECT 364.995 -2.205 365.325 -1.875 ;
        RECT 363.635 -2.205 363.965 -1.875 ;
        RECT 362.275 -2.205 362.605 -1.875 ;
        RECT 360.915 -2.205 361.245 -1.875 ;
        RECT 359.555 -2.205 359.885 -1.875 ;
        RECT 358.195 -2.205 358.525 -1.875 ;
        RECT 356.835 -2.205 357.165 -1.875 ;
        RECT 355.475 -2.205 355.805 -1.875 ;
        RECT 354.115 -2.205 354.445 -1.875 ;
        RECT 352.755 -2.205 353.085 -1.875 ;
        RECT 351.395 -2.205 351.725 -1.875 ;
        RECT 350.035 -2.205 350.365 -1.875 ;
        RECT 348.675 -2.205 349.005 -1.875 ;
        RECT 347.315 -2.205 347.645 -1.875 ;
        RECT 345.955 -2.205 346.285 -1.875 ;
        RECT 344.595 -2.205 344.925 -1.875 ;
        RECT 343.235 -2.205 343.565 -1.875 ;
        RECT 341.875 -2.205 342.205 -1.875 ;
        RECT 340.515 -2.205 340.845 -1.875 ;
        RECT 339.155 -2.205 339.485 -1.875 ;
        RECT 337.795 -2.205 338.125 -1.875 ;
        RECT 336.435 -2.205 336.765 -1.875 ;
        RECT 335.075 -2.205 335.405 -1.875 ;
        RECT 333.715 -2.205 334.045 -1.875 ;
        RECT 332.355 -2.205 332.685 -1.875 ;
        RECT 330.995 -2.205 331.325 -1.875 ;
        RECT 329.635 -2.205 329.965 -1.875 ;
        RECT 328.275 -2.205 328.605 -1.875 ;
        RECT 326.915 -2.205 327.245 -1.875 ;
        RECT 325.555 -2.205 325.885 -1.875 ;
        RECT 324.195 -2.205 324.525 -1.875 ;
        RECT 322.835 -2.205 323.165 -1.875 ;
        RECT 321.475 -2.205 321.805 -1.875 ;
        RECT 320.115 -2.205 320.445 -1.875 ;
        RECT 318.755 -2.205 319.085 -1.875 ;
        RECT 317.395 -2.205 317.725 -1.875 ;
        RECT 316.035 -2.205 316.365 -1.875 ;
        RECT 314.675 -2.205 315.005 -1.875 ;
        RECT 313.315 -2.205 313.645 -1.875 ;
        RECT 311.955 -2.205 312.285 -1.875 ;
        RECT 310.595 -2.205 310.925 -1.875 ;
        RECT 309.235 -2.205 309.565 -1.875 ;
        RECT 307.875 -2.205 308.205 -1.875 ;
        RECT 306.515 -2.205 306.845 -1.875 ;
        RECT 305.155 -2.205 305.485 -1.875 ;
        RECT 303.795 -2.205 304.125 -1.875 ;
        RECT 302.435 -2.205 302.765 -1.875 ;
        RECT 301.075 -2.205 301.405 -1.875 ;
        RECT 299.715 -2.205 300.045 -1.875 ;
        RECT 298.355 -2.205 298.685 -1.875 ;
        RECT 296.995 -2.205 297.325 -1.875 ;
        RECT 295.635 -2.205 295.965 -1.875 ;
        RECT 294.275 -2.205 294.605 -1.875 ;
        RECT 292.915 -2.205 293.245 -1.875 ;
        RECT 291.555 -2.205 291.885 -1.875 ;
        RECT 290.195 -2.205 290.525 -1.875 ;
        RECT 288.835 -2.205 289.165 -1.875 ;
        RECT 287.475 -2.205 287.805 -1.875 ;
        RECT 286.115 -2.205 286.445 -1.875 ;
        RECT 284.755 -2.205 285.085 -1.875 ;
        RECT 283.395 -2.205 283.725 -1.875 ;
        RECT 282.035 -2.205 282.365 -1.875 ;
        RECT 280.675 -2.205 281.005 -1.875 ;
        RECT 279.315 -2.205 279.645 -1.875 ;
        RECT 277.955 -2.205 278.285 -1.875 ;
        RECT 276.595 -2.205 276.925 -1.875 ;
        RECT 275.235 -2.205 275.565 -1.875 ;
        RECT 273.875 -2.205 274.205 -1.875 ;
        RECT 272.515 -2.205 272.845 -1.875 ;
        RECT 271.155 -2.205 271.485 -1.875 ;
        RECT 269.795 -2.205 270.125 -1.875 ;
        RECT 268.435 -2.205 268.765 -1.875 ;
        RECT 267.075 -2.205 267.405 -1.875 ;
        RECT 265.715 -2.205 266.045 -1.875 ;
        RECT 264.355 -2.205 264.685 -1.875 ;
        RECT 262.995 -2.205 263.325 -1.875 ;
        RECT 261.635 -2.205 261.965 -1.875 ;
        RECT 260.275 -2.205 260.605 -1.875 ;
        RECT 258.915 -2.205 259.245 -1.875 ;
        RECT 257.555 -2.205 257.885 -1.875 ;
        RECT 256.195 -2.205 256.525 -1.875 ;
        RECT 254.835 -2.205 255.165 -1.875 ;
        RECT 253.475 -2.205 253.805 -1.875 ;
        RECT 252.115 -2.205 252.445 -1.875 ;
        RECT 250.755 -2.205 251.085 -1.875 ;
        RECT 249.395 -2.205 249.725 -1.875 ;
        RECT 248.035 -2.205 248.365 -1.875 ;
        RECT 246.675 -2.205 247.005 -1.875 ;
        RECT 245.315 -2.205 245.645 -1.875 ;
        RECT 243.955 -2.205 244.285 -1.875 ;
        RECT 242.595 -2.205 242.925 -1.875 ;
        RECT 241.235 -2.205 241.565 -1.875 ;
        RECT 239.875 -2.205 240.205 -1.875 ;
        RECT 238.515 -2.205 238.845 -1.875 ;
        RECT 237.155 -2.205 237.485 -1.875 ;
        RECT 235.795 -2.205 236.125 -1.875 ;
        RECT 234.435 -2.205 234.765 -1.875 ;
        RECT 233.075 -2.205 233.405 -1.875 ;
        RECT 231.715 -2.205 232.045 -1.875 ;
        RECT 230.355 -2.205 230.685 -1.875 ;
        RECT 228.995 -2.205 229.325 -1.875 ;
        RECT 227.635 -2.205 227.965 -1.875 ;
        RECT 226.275 -2.205 226.605 -1.875 ;
        RECT 224.915 -2.205 225.245 -1.875 ;
        RECT 223.555 -2.205 223.885 -1.875 ;
        RECT 222.195 -2.205 222.525 -1.875 ;
        RECT 220.835 -2.205 221.165 -1.875 ;
        RECT 219.475 -2.205 219.805 -1.875 ;
        RECT 218.115 -2.205 218.445 -1.875 ;
        RECT 216.755 -2.205 217.085 -1.875 ;
        RECT 215.395 -2.205 215.725 -1.875 ;
        RECT 214.035 -2.205 214.365 -1.875 ;
        RECT 212.675 -2.205 213.005 -1.875 ;
        RECT 211.315 -2.205 211.645 -1.875 ;
        RECT 209.955 -2.205 210.285 -1.875 ;
        RECT 208.595 -2.205 208.925 -1.875 ;
        RECT 207.235 -2.205 207.565 -1.875 ;
        RECT 205.875 -2.205 206.205 -1.875 ;
        RECT 204.515 -2.205 204.845 -1.875 ;
        RECT 203.155 -2.205 203.485 -1.875 ;
        RECT 201.795 -2.205 202.125 -1.875 ;
        RECT 200.435 -2.205 200.765 -1.875 ;
        RECT 199.075 -2.205 199.405 -1.875 ;
        RECT 197.715 -2.205 198.045 -1.875 ;
        RECT 196.355 -2.205 196.685 -1.875 ;
        RECT 194.995 -2.205 195.325 -1.875 ;
        RECT 193.635 -2.205 193.965 -1.875 ;
        RECT 192.275 -2.205 192.605 -1.875 ;
        RECT 190.915 -2.205 191.245 -1.875 ;
        RECT 189.555 -2.205 189.885 -1.875 ;
        RECT 188.195 -2.205 188.525 -1.875 ;
        RECT 186.835 -2.205 187.165 -1.875 ;
        RECT 185.475 -2.205 185.805 -1.875 ;
        RECT 184.115 -2.205 184.445 -1.875 ;
        RECT 182.755 -2.205 183.085 -1.875 ;
        RECT 181.395 -2.205 181.725 -1.875 ;
        RECT 180.035 -2.205 180.365 -1.875 ;
        RECT 178.675 -2.205 179.005 -1.875 ;
        RECT 177.315 -2.205 177.645 -1.875 ;
        RECT 175.955 -2.205 176.285 -1.875 ;
        RECT 174.595 -2.205 174.925 -1.875 ;
        RECT 173.235 -2.205 173.565 -1.875 ;
        RECT 171.875 -2.205 172.205 -1.875 ;
        RECT 170.515 -2.205 170.845 -1.875 ;
        RECT 169.155 -2.205 169.485 -1.875 ;
        RECT 167.795 -2.205 168.125 -1.875 ;
        RECT 166.435 -2.205 166.765 -1.875 ;
        RECT 165.075 -2.205 165.405 -1.875 ;
        RECT 163.715 -2.205 164.045 -1.875 ;
        RECT 162.355 -2.205 162.685 -1.875 ;
        RECT 160.995 -2.205 161.325 -1.875 ;
        RECT 159.635 -2.205 159.965 -1.875 ;
        RECT 158.275 -2.205 158.605 -1.875 ;
        RECT 156.915 -2.205 157.245 -1.875 ;
        RECT 155.555 -2.205 155.885 -1.875 ;
        RECT 154.195 -2.205 154.525 -1.875 ;
        RECT 152.835 -2.205 153.165 -1.875 ;
        RECT 151.475 -2.205 151.805 -1.875 ;
        RECT 150.115 -2.205 150.445 -1.875 ;
        RECT 148.755 -2.205 149.085 -1.875 ;
        RECT 147.395 -2.205 147.725 -1.875 ;
        RECT 146.035 -2.205 146.365 -1.875 ;
        RECT 144.675 -2.205 145.005 -1.875 ;
        RECT 143.315 -2.205 143.645 -1.875 ;
        RECT 141.955 -2.205 142.285 -1.875 ;
        RECT 140.595 -2.205 140.925 -1.875 ;
        RECT 139.235 -2.205 139.565 -1.875 ;
        RECT 137.875 -2.205 138.205 -1.875 ;
        RECT 136.515 -2.205 136.845 -1.875 ;
        RECT 135.155 -2.205 135.485 -1.875 ;
        RECT 133.795 -2.205 134.125 -1.875 ;
        RECT 132.435 -2.205 132.765 -1.875 ;
        RECT 131.075 -2.205 131.405 -1.875 ;
        RECT 129.715 -2.205 130.045 -1.875 ;
        RECT 128.355 -2.205 128.685 -1.875 ;
        RECT 126.995 -2.205 127.325 -1.875 ;
        RECT 125.635 -2.205 125.965 -1.875 ;
        RECT 124.275 -2.205 124.605 -1.875 ;
        RECT 122.915 -2.205 123.245 -1.875 ;
        RECT 121.555 -2.205 121.885 -1.875 ;
        RECT 120.195 -2.205 120.525 -1.875 ;
        RECT 118.835 -2.205 119.165 -1.875 ;
        RECT 117.475 -2.205 117.805 -1.875 ;
        RECT 116.115 -2.205 116.445 -1.875 ;
        RECT 114.755 -2.205 115.085 -1.875 ;
        RECT 113.395 -2.205 113.725 -1.875 ;
        RECT 112.035 -2.205 112.365 -1.875 ;
        RECT 110.675 -2.205 111.005 -1.875 ;
        RECT 109.315 -2.205 109.645 -1.875 ;
        RECT 107.955 -2.205 108.285 -1.875 ;
        RECT 106.595 -2.205 106.925 -1.875 ;
        RECT 105.235 -2.205 105.565 -1.875 ;
        RECT 103.875 -2.205 104.205 -1.875 ;
        RECT 102.515 -2.205 102.845 -1.875 ;
        RECT 101.155 -2.205 101.485 -1.875 ;
        RECT 99.795 -2.205 100.125 -1.875 ;
        RECT 98.435 -2.205 98.765 -1.875 ;
        RECT 97.075 -2.205 97.405 -1.875 ;
        RECT 95.715 -2.205 96.045 -1.875 ;
        RECT 94.355 -2.205 94.685 -1.875 ;
        RECT 92.995 -2.205 93.325 -1.875 ;
        RECT 91.635 -2.205 91.965 -1.875 ;
        RECT 90.275 -2.205 90.605 -1.875 ;
        RECT 88.915 -2.205 89.245 -1.875 ;
        RECT 87.555 -2.205 87.885 -1.875 ;
        RECT 86.195 -2.205 86.525 -1.875 ;
        RECT 84.835 -2.205 85.165 -1.875 ;
        RECT 83.475 -2.205 83.805 -1.875 ;
        RECT 82.115 -2.205 82.445 -1.875 ;
        RECT 80.755 -2.205 81.085 -1.875 ;
        RECT 79.395 -2.205 79.725 -1.875 ;
        RECT 78.035 -2.205 78.365 -1.875 ;
        RECT 76.675 -2.205 77.005 -1.875 ;
        RECT 75.315 -2.205 75.645 -1.875 ;
        RECT 73.955 -2.205 74.285 -1.875 ;
        RECT 72.595 -2.205 72.925 -1.875 ;
        RECT 71.235 -2.205 71.565 -1.875 ;
        RECT 69.875 -2.205 70.205 -1.875 ;
        RECT 68.515 -2.205 68.845 -1.875 ;
        RECT 67.155 -2.205 67.485 -1.875 ;
        RECT 65.795 -2.205 66.125 -1.875 ;
        RECT 64.435 -2.205 64.765 -1.875 ;
        RECT 63.075 -2.205 63.405 -1.875 ;
        RECT 61.715 -2.205 62.045 -1.875 ;
        RECT 60.355 -2.205 60.685 -1.875 ;
        RECT 58.995 -2.205 59.325 -1.875 ;
        RECT 57.635 -2.205 57.965 -1.875 ;
        RECT 56.275 -2.205 56.605 -1.875 ;
        RECT 54.915 -2.205 55.245 -1.875 ;
        RECT 53.555 -2.205 53.885 -1.875 ;
        RECT 52.195 -2.205 52.525 -1.875 ;
        RECT 50.835 -2.205 51.165 -1.875 ;
        RECT 49.475 -2.205 49.805 -1.875 ;
        RECT 48.115 -2.205 48.445 -1.875 ;
        RECT 46.755 -2.205 47.085 -1.875 ;
        RECT 45.395 -2.205 45.725 -1.875 ;
        RECT 44.035 -2.205 44.365 -1.875 ;
        RECT 42.675 -2.205 43.005 -1.875 ;
        RECT 41.315 -2.205 41.645 -1.875 ;
        RECT 39.955 -2.205 40.285 -1.875 ;
        RECT 38.595 -2.205 38.925 -1.875 ;
        RECT 37.235 -2.205 37.565 -1.875 ;
        RECT 35.875 -2.205 36.205 -1.875 ;
        RECT 34.515 -2.205 34.845 -1.875 ;
        RECT 33.155 -2.205 33.485 -1.875 ;
        RECT 31.795 -2.205 32.125 -1.875 ;
        RECT 30.435 -2.205 30.765 -1.875 ;
        RECT 29.075 -2.205 29.405 -1.875 ;
        RECT 27.715 -2.205 28.045 -1.875 ;
        RECT 26.355 -2.205 26.685 -1.875 ;
        RECT 24.995 -2.205 25.325 -1.875 ;
        RECT 23.635 -2.205 23.965 -1.875 ;
        RECT 22.275 -2.205 22.605 -1.875 ;
        RECT 20.915 -2.205 21.245 -1.875 ;
        RECT 19.555 -2.205 19.885 -1.875 ;
        RECT 18.195 -2.205 18.525 -1.875 ;
        RECT 16.835 -2.205 17.165 -1.875 ;
        RECT 15.475 -2.205 15.805 -1.875 ;
        RECT 14.115 -2.205 14.445 -1.875 ;
        RECT 12.755 -2.205 13.085 -1.875 ;
        RECT 11.395 -2.205 11.725 -1.875 ;
        RECT 10.035 -2.205 10.365 -1.875 ;
        RECT 8.675 -2.205 9.005 -1.875 ;
        RECT 7.315 -2.205 7.645 -1.875 ;
        RECT 5.955 -2.205 6.285 -1.875 ;
        RECT 4.595 -2.205 4.925 -1.875 ;
        RECT 3.235 -2.205 3.565 -1.875 ;
        RECT 1.875 -2.205 2.205 -1.875 ;
        RECT 0.515 -2.205 0.845 -1.875 ;
        RECT -0.845 -2.205 -0.515 -1.875 ;
        RECT 678.125 -2.2 954.88 -1.88 ;
        RECT 953.875 -2.205 954.205 -1.875 ;
        RECT 952.515 -2.205 952.845 -1.875 ;
        RECT 951.155 -2.205 951.485 -1.875 ;
        RECT 949.795 -2.205 950.125 -1.875 ;
        RECT 948.435 -2.205 948.765 -1.875 ;
        RECT 947.075 -2.205 947.405 -1.875 ;
        RECT 945.715 -2.205 946.045 -1.875 ;
        RECT 944.355 -2.205 944.685 -1.875 ;
        RECT 942.995 -2.205 943.325 -1.875 ;
        RECT 941.635 -2.205 941.965 -1.875 ;
        RECT 940.275 -2.205 940.605 -1.875 ;
        RECT 938.915 -2.205 939.245 -1.875 ;
        RECT 937.555 -2.205 937.885 -1.875 ;
        RECT 936.195 -2.205 936.525 -1.875 ;
        RECT 934.835 -2.205 935.165 -1.875 ;
        RECT 933.475 -2.205 933.805 -1.875 ;
        RECT 932.115 -2.205 932.445 -1.875 ;
        RECT 930.755 -2.205 931.085 -1.875 ;
        RECT 929.395 -2.205 929.725 -1.875 ;
        RECT 928.035 -2.205 928.365 -1.875 ;
        RECT 926.675 -2.205 927.005 -1.875 ;
        RECT 925.315 -2.205 925.645 -1.875 ;
        RECT 923.955 -2.205 924.285 -1.875 ;
        RECT 922.595 -2.205 922.925 -1.875 ;
        RECT 921.235 -2.205 921.565 -1.875 ;
        RECT 919.875 -2.205 920.205 -1.875 ;
        RECT 918.515 -2.205 918.845 -1.875 ;
        RECT 917.155 -2.205 917.485 -1.875 ;
        RECT 915.795 -2.205 916.125 -1.875 ;
        RECT 914.435 -2.205 914.765 -1.875 ;
        RECT 913.075 -2.205 913.405 -1.875 ;
        RECT 911.715 -2.205 912.045 -1.875 ;
        RECT 910.355 -2.205 910.685 -1.875 ;
        RECT 908.995 -2.205 909.325 -1.875 ;
        RECT 907.635 -2.205 907.965 -1.875 ;
        RECT 906.275 -2.205 906.605 -1.875 ;
        RECT 904.915 -2.205 905.245 -1.875 ;
        RECT 903.555 -2.205 903.885 -1.875 ;
        RECT 902.195 -2.205 902.525 -1.875 ;
        RECT 900.835 -2.205 901.165 -1.875 ;
        RECT 899.475 -2.205 899.805 -1.875 ;
        RECT 898.115 -2.205 898.445 -1.875 ;
        RECT 896.755 -2.205 897.085 -1.875 ;
        RECT 895.395 -2.205 895.725 -1.875 ;
        RECT 894.035 -2.205 894.365 -1.875 ;
        RECT 892.675 -2.205 893.005 -1.875 ;
        RECT 891.315 -2.205 891.645 -1.875 ;
        RECT 889.955 -2.205 890.285 -1.875 ;
        RECT 888.595 -2.205 888.925 -1.875 ;
        RECT 887.235 -2.205 887.565 -1.875 ;
        RECT 885.875 -2.205 886.205 -1.875 ;
        RECT 884.515 -2.205 884.845 -1.875 ;
        RECT 883.155 -2.205 883.485 -1.875 ;
        RECT 881.795 -2.205 882.125 -1.875 ;
        RECT 880.435 -2.205 880.765 -1.875 ;
        RECT 879.075 -2.205 879.405 -1.875 ;
        RECT 877.715 -2.205 878.045 -1.875 ;
        RECT 876.355 -2.205 876.685 -1.875 ;
        RECT 874.995 -2.205 875.325 -1.875 ;
        RECT 873.635 -2.205 873.965 -1.875 ;
        RECT 872.275 -2.205 872.605 -1.875 ;
        RECT 870.915 -2.205 871.245 -1.875 ;
        RECT 869.555 -2.205 869.885 -1.875 ;
        RECT 868.195 -2.205 868.525 -1.875 ;
        RECT 866.835 -2.205 867.165 -1.875 ;
        RECT 865.475 -2.205 865.805 -1.875 ;
        RECT 864.115 -2.205 864.445 -1.875 ;
        RECT 862.755 -2.205 863.085 -1.875 ;
        RECT 861.395 -2.205 861.725 -1.875 ;
        RECT 860.035 -2.205 860.365 -1.875 ;
        RECT 858.675 -2.205 859.005 -1.875 ;
        RECT 857.315 -2.205 857.645 -1.875 ;
        RECT 855.955 -2.205 856.285 -1.875 ;
        RECT 854.595 -2.205 854.925 -1.875 ;
        RECT 853.235 -2.205 853.565 -1.875 ;
        RECT 851.875 -2.205 852.205 -1.875 ;
        RECT 850.515 -2.205 850.845 -1.875 ;
        RECT 849.155 -2.205 849.485 -1.875 ;
        RECT 847.795 -2.205 848.125 -1.875 ;
        RECT 846.435 -2.205 846.765 -1.875 ;
        RECT 845.075 -2.205 845.405 -1.875 ;
        RECT 843.715 -2.205 844.045 -1.875 ;
        RECT 842.355 -2.205 842.685 -1.875 ;
        RECT 840.995 -2.205 841.325 -1.875 ;
        RECT 839.635 -2.205 839.965 -1.875 ;
        RECT 838.275 -2.205 838.605 -1.875 ;
        RECT 836.915 -2.205 837.245 -1.875 ;
        RECT 835.555 -2.205 835.885 -1.875 ;
        RECT 834.195 -2.205 834.525 -1.875 ;
        RECT 832.835 -2.205 833.165 -1.875 ;
        RECT 831.475 -2.205 831.805 -1.875 ;
        RECT 830.115 -2.205 830.445 -1.875 ;
        RECT 828.755 -2.205 829.085 -1.875 ;
        RECT 827.395 -2.205 827.725 -1.875 ;
        RECT 826.035 -2.205 826.365 -1.875 ;
        RECT 824.675 -2.205 825.005 -1.875 ;
        RECT 823.315 -2.205 823.645 -1.875 ;
        RECT 821.955 -2.205 822.285 -1.875 ;
        RECT 820.595 -2.205 820.925 -1.875 ;
        RECT 819.235 -2.205 819.565 -1.875 ;
        RECT 817.875 -2.205 818.205 -1.875 ;
        RECT 816.515 -2.205 816.845 -1.875 ;
        RECT 815.155 -2.205 815.485 -1.875 ;
        RECT 813.795 -2.205 814.125 -1.875 ;
        RECT 812.435 -2.205 812.765 -1.875 ;
        RECT 811.075 -2.205 811.405 -1.875 ;
        RECT 809.715 -2.205 810.045 -1.875 ;
        RECT 808.355 -2.205 808.685 -1.875 ;
        RECT 806.995 -2.205 807.325 -1.875 ;
        RECT 805.635 -2.205 805.965 -1.875 ;
        RECT 804.275 -2.205 804.605 -1.875 ;
        RECT 802.915 -2.205 803.245 -1.875 ;
        RECT 801.555 -2.205 801.885 -1.875 ;
        RECT 800.195 -2.205 800.525 -1.875 ;
        RECT 798.835 -2.205 799.165 -1.875 ;
        RECT 797.475 -2.205 797.805 -1.875 ;
        RECT 796.115 -2.205 796.445 -1.875 ;
        RECT 794.755 -2.205 795.085 -1.875 ;
        RECT 793.395 -2.205 793.725 -1.875 ;
        RECT 792.035 -2.205 792.365 -1.875 ;
        RECT 790.675 -2.205 791.005 -1.875 ;
        RECT 789.315 -2.205 789.645 -1.875 ;
        RECT 787.955 -2.205 788.285 -1.875 ;
        RECT 786.595 -2.205 786.925 -1.875 ;
        RECT 785.235 -2.205 785.565 -1.875 ;
        RECT 783.875 -2.205 784.205 -1.875 ;
        RECT 782.515 -2.205 782.845 -1.875 ;
        RECT 781.155 -2.205 781.485 -1.875 ;
        RECT 779.795 -2.205 780.125 -1.875 ;
        RECT 778.435 -2.205 778.765 -1.875 ;
        RECT 777.075 -2.205 777.405 -1.875 ;
        RECT 775.715 -2.205 776.045 -1.875 ;
        RECT 774.355 -2.205 774.685 -1.875 ;
        RECT 772.995 -2.205 773.325 -1.875 ;
        RECT 771.635 -2.205 771.965 -1.875 ;
        RECT 770.275 -2.205 770.605 -1.875 ;
        RECT 768.915 -2.205 769.245 -1.875 ;
        RECT 767.555 -2.205 767.885 -1.875 ;
        RECT 766.195 -2.205 766.525 -1.875 ;
        RECT 764.835 -2.205 765.165 -1.875 ;
        RECT 763.475 -2.205 763.805 -1.875 ;
        RECT 762.115 -2.205 762.445 -1.875 ;
        RECT 760.755 -2.205 761.085 -1.875 ;
        RECT 759.395 -2.205 759.725 -1.875 ;
        RECT 758.035 -2.205 758.365 -1.875 ;
        RECT 756.675 -2.205 757.005 -1.875 ;
        RECT 755.315 -2.205 755.645 -1.875 ;
        RECT 753.955 -2.205 754.285 -1.875 ;
        RECT 752.595 -2.205 752.925 -1.875 ;
        RECT 751.235 -2.205 751.565 -1.875 ;
        RECT 749.875 -2.205 750.205 -1.875 ;
        RECT 748.515 -2.205 748.845 -1.875 ;
        RECT 747.155 -2.205 747.485 -1.875 ;
        RECT 745.795 -2.205 746.125 -1.875 ;
        RECT 744.435 -2.205 744.765 -1.875 ;
        RECT 743.075 -2.205 743.405 -1.875 ;
        RECT 741.715 -2.205 742.045 -1.875 ;
        RECT 740.355 -2.205 740.685 -1.875 ;
        RECT 738.995 -2.205 739.325 -1.875 ;
        RECT 737.635 -2.205 737.965 -1.875 ;
        RECT 736.275 -2.205 736.605 -1.875 ;
        RECT 734.915 -2.205 735.245 -1.875 ;
        RECT 733.555 -2.205 733.885 -1.875 ;
        RECT 732.195 -2.205 732.525 -1.875 ;
        RECT 730.835 -2.205 731.165 -1.875 ;
        RECT 729.475 -2.205 729.805 -1.875 ;
        RECT 728.115 -2.205 728.445 -1.875 ;
        RECT 726.755 -2.205 727.085 -1.875 ;
        RECT 725.395 -2.205 725.725 -1.875 ;
        RECT 724.035 -2.205 724.365 -1.875 ;
        RECT 722.675 -2.205 723.005 -1.875 ;
        RECT 721.315 -2.205 721.645 -1.875 ;
        RECT 719.955 -2.205 720.285 -1.875 ;
        RECT 718.595 -2.205 718.925 -1.875 ;
        RECT 717.235 -2.205 717.565 -1.875 ;
        RECT 715.875 -2.205 716.205 -1.875 ;
        RECT 714.515 -2.205 714.845 -1.875 ;
        RECT 713.155 -2.205 713.485 -1.875 ;
        RECT 711.795 -2.205 712.125 -1.875 ;
        RECT 710.435 -2.205 710.765 -1.875 ;
        RECT 709.075 -2.205 709.405 -1.875 ;
        RECT 707.715 -2.205 708.045 -1.875 ;
        RECT 706.355 -2.205 706.685 -1.875 ;
        RECT 704.995 -2.205 705.325 -1.875 ;
        RECT 703.635 -2.205 703.965 -1.875 ;
        RECT 702.275 -2.205 702.605 -1.875 ;
        RECT 700.915 -2.205 701.245 -1.875 ;
        RECT 699.555 -2.205 699.885 -1.875 ;
        RECT 698.195 -2.205 698.525 -1.875 ;
        RECT 696.835 -2.205 697.165 -1.875 ;
        RECT 695.475 -2.205 695.805 -1.875 ;
        RECT 694.115 -2.205 694.445 -1.875 ;
        RECT 692.755 -2.205 693.085 -1.875 ;
        RECT 691.395 -2.205 691.725 -1.875 ;
        RECT 690.035 -2.205 690.365 -1.875 ;
        RECT 688.675 -2.205 689.005 -1.875 ;
        RECT 687.315 -2.205 687.645 -1.875 ;
        RECT 685.955 -2.205 686.285 -1.875 ;
        RECT 684.595 -2.205 684.925 -1.875 ;
        RECT 683.235 -2.205 683.565 -1.875 ;
        RECT 681.875 -2.205 682.205 -1.875 ;
        RECT 680.515 -2.205 680.845 -1.875 ;
        RECT 679.155 -2.205 679.485 -1.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -3.565 136.845 -3.235 ;
        RECT 135.155 -3.565 135.485 -3.235 ;
        RECT 133.795 -3.565 134.125 -3.235 ;
        RECT 132.435 -3.565 132.765 -3.235 ;
        RECT 131.075 -3.565 131.405 -3.235 ;
        RECT 129.715 -3.565 130.045 -3.235 ;
        RECT 128.355 -3.565 128.685 -3.235 ;
        RECT 126.995 -3.565 127.325 -3.235 ;
        RECT 125.635 -3.565 125.965 -3.235 ;
        RECT 124.275 -3.565 124.605 -3.235 ;
        RECT 122.915 -3.565 123.245 -3.235 ;
        RECT 121.555 -3.565 121.885 -3.235 ;
        RECT 120.195 -3.565 120.525 -3.235 ;
        RECT 118.835 -3.565 119.165 -3.235 ;
        RECT 117.475 -3.565 117.805 -3.235 ;
        RECT 116.115 -3.565 116.445 -3.235 ;
        RECT 114.755 -3.565 115.085 -3.235 ;
        RECT 113.395 -3.565 113.725 -3.235 ;
        RECT 112.035 -3.565 112.365 -3.235 ;
        RECT 110.675 -3.565 111.005 -3.235 ;
        RECT 109.315 -3.565 109.645 -3.235 ;
        RECT 107.955 -3.565 108.285 -3.235 ;
        RECT 106.595 -3.565 106.925 -3.235 ;
        RECT 105.235 -3.565 105.565 -3.235 ;
        RECT 103.875 -3.565 104.205 -3.235 ;
        RECT 102.515 -3.565 102.845 -3.235 ;
        RECT 101.155 -3.565 101.485 -3.235 ;
        RECT 99.795 -3.565 100.125 -3.235 ;
        RECT 98.435 -3.565 98.765 -3.235 ;
        RECT 97.075 -3.565 97.405 -3.235 ;
        RECT 95.715 -3.565 96.045 -3.235 ;
        RECT 94.355 -3.565 94.685 -3.235 ;
        RECT 92.995 -3.565 93.325 -3.235 ;
        RECT 91.635 -3.565 91.965 -3.235 ;
        RECT 90.275 -3.565 90.605 -3.235 ;
        RECT 88.915 -3.565 89.245 -3.235 ;
        RECT 87.555 -3.565 87.885 -3.235 ;
        RECT 86.195 -3.565 86.525 -3.235 ;
        RECT 84.835 -3.565 85.165 -3.235 ;
        RECT 83.475 -3.565 83.805 -3.235 ;
        RECT 82.115 -3.565 82.445 -3.235 ;
        RECT 80.755 -3.565 81.085 -3.235 ;
        RECT 79.395 -3.565 79.725 -3.235 ;
        RECT 78.035 -3.565 78.365 -3.235 ;
        RECT 76.675 -3.565 77.005 -3.235 ;
        RECT 75.315 -3.565 75.645 -3.235 ;
        RECT 73.955 -3.565 74.285 -3.235 ;
        RECT 72.595 -3.565 72.925 -3.235 ;
        RECT 71.235 -3.565 71.565 -3.235 ;
        RECT 69.875 -3.565 70.205 -3.235 ;
        RECT 68.515 -3.565 68.845 -3.235 ;
        RECT 67.155 -3.565 67.485 -3.235 ;
        RECT 65.795 -3.565 66.125 -3.235 ;
        RECT 64.435 -3.565 64.765 -3.235 ;
        RECT 63.075 -3.565 63.405 -3.235 ;
        RECT 61.715 -3.565 62.045 -3.235 ;
        RECT 60.355 -3.565 60.685 -3.235 ;
        RECT 58.995 -3.565 59.325 -3.235 ;
        RECT 57.635 -3.565 57.965 -3.235 ;
        RECT 56.275 -3.565 56.605 -3.235 ;
        RECT 54.915 -3.565 55.245 -3.235 ;
        RECT 53.555 -3.565 53.885 -3.235 ;
        RECT 52.195 -3.565 52.525 -3.235 ;
        RECT 50.835 -3.565 51.165 -3.235 ;
        RECT 49.475 -3.565 49.805 -3.235 ;
        RECT 48.115 -3.565 48.445 -3.235 ;
        RECT 46.755 -3.565 47.085 -3.235 ;
        RECT 45.395 -3.565 45.725 -3.235 ;
        RECT 44.035 -3.565 44.365 -3.235 ;
        RECT 42.675 -3.565 43.005 -3.235 ;
        RECT 41.315 -3.565 41.645 -3.235 ;
        RECT 39.955 -3.565 40.285 -3.235 ;
        RECT 38.595 -3.565 38.925 -3.235 ;
        RECT 37.235 -3.565 37.565 -3.235 ;
        RECT 35.875 -3.565 36.205 -3.235 ;
        RECT 34.515 -3.565 34.845 -3.235 ;
        RECT 33.155 -3.565 33.485 -3.235 ;
        RECT 31.795 -3.565 32.125 -3.235 ;
        RECT 30.435 -3.565 30.765 -3.235 ;
        RECT 29.075 -3.565 29.405 -3.235 ;
        RECT 27.715 -3.565 28.045 -3.235 ;
        RECT 26.355 -3.565 26.685 -3.235 ;
        RECT 24.995 -3.565 25.325 -3.235 ;
        RECT 23.635 -3.565 23.965 -3.235 ;
        RECT 22.275 -3.565 22.605 -3.235 ;
        RECT 20.915 -3.565 21.245 -3.235 ;
        RECT 19.555 -3.565 19.885 -3.235 ;
        RECT 18.195 -3.565 18.525 -3.235 ;
        RECT 16.835 -3.565 17.165 -3.235 ;
        RECT 15.475 -3.565 15.805 -3.235 ;
        RECT 14.115 -3.565 14.445 -3.235 ;
        RECT 12.755 -3.565 13.085 -3.235 ;
        RECT 11.395 -3.565 11.725 -3.235 ;
        RECT 10.035 -3.565 10.365 -3.235 ;
        RECT 8.675 -3.565 9.005 -3.235 ;
        RECT 7.315 -3.565 7.645 -3.235 ;
        RECT 5.955 -3.565 6.285 -3.235 ;
        RECT 4.595 -3.565 4.925 -3.235 ;
        RECT 3.235 -3.565 3.565 -3.235 ;
        RECT 1.875 -3.565 2.205 -3.235 ;
        RECT 0.515 -3.565 0.845 -3.235 ;
        RECT -0.845 -3.565 -0.515 -3.235 ;
        RECT 677.795 -3.565 678.125 -3.235 ;
        RECT -1.52 -3.56 678.125 -3.24 ;
        RECT 676.435 -3.565 676.765 -3.235 ;
        RECT 675.075 -3.565 675.405 -3.235 ;
        RECT 673.715 -3.565 674.045 -3.235 ;
        RECT 672.355 -3.565 672.685 -3.235 ;
        RECT 670.995 -3.565 671.325 -3.235 ;
        RECT 669.635 -3.565 669.965 -3.235 ;
        RECT 668.275 -3.565 668.605 -3.235 ;
        RECT 666.915 -3.565 667.245 -3.235 ;
        RECT 665.555 -3.565 665.885 -3.235 ;
        RECT 664.195 -3.565 664.525 -3.235 ;
        RECT 662.835 -3.565 663.165 -3.235 ;
        RECT 661.475 -3.565 661.805 -3.235 ;
        RECT 660.115 -3.565 660.445 -3.235 ;
        RECT 658.755 -3.565 659.085 -3.235 ;
        RECT 657.395 -3.565 657.725 -3.235 ;
        RECT 656.035 -3.565 656.365 -3.235 ;
        RECT 654.675 -3.565 655.005 -3.235 ;
        RECT 653.315 -3.565 653.645 -3.235 ;
        RECT 651.955 -3.565 652.285 -3.235 ;
        RECT 650.595 -3.565 650.925 -3.235 ;
        RECT 649.235 -3.565 649.565 -3.235 ;
        RECT 647.875 -3.565 648.205 -3.235 ;
        RECT 646.515 -3.565 646.845 -3.235 ;
        RECT 645.155 -3.565 645.485 -3.235 ;
        RECT 643.795 -3.565 644.125 -3.235 ;
        RECT 642.435 -3.565 642.765 -3.235 ;
        RECT 641.075 -3.565 641.405 -3.235 ;
        RECT 639.715 -3.565 640.045 -3.235 ;
        RECT 638.355 -3.565 638.685 -3.235 ;
        RECT 636.995 -3.565 637.325 -3.235 ;
        RECT 635.635 -3.565 635.965 -3.235 ;
        RECT 634.275 -3.565 634.605 -3.235 ;
        RECT 632.915 -3.565 633.245 -3.235 ;
        RECT 631.555 -3.565 631.885 -3.235 ;
        RECT 630.195 -3.565 630.525 -3.235 ;
        RECT 628.835 -3.565 629.165 -3.235 ;
        RECT 627.475 -3.565 627.805 -3.235 ;
        RECT 626.115 -3.565 626.445 -3.235 ;
        RECT 624.755 -3.565 625.085 -3.235 ;
        RECT 623.395 -3.565 623.725 -3.235 ;
        RECT 622.035 -3.565 622.365 -3.235 ;
        RECT 620.675 -3.565 621.005 -3.235 ;
        RECT 619.315 -3.565 619.645 -3.235 ;
        RECT 617.955 -3.565 618.285 -3.235 ;
        RECT 616.595 -3.565 616.925 -3.235 ;
        RECT 615.235 -3.565 615.565 -3.235 ;
        RECT 613.875 -3.565 614.205 -3.235 ;
        RECT 612.515 -3.565 612.845 -3.235 ;
        RECT 611.155 -3.565 611.485 -3.235 ;
        RECT 609.795 -3.565 610.125 -3.235 ;
        RECT 608.435 -3.565 608.765 -3.235 ;
        RECT 607.075 -3.565 607.405 -3.235 ;
        RECT 605.715 -3.565 606.045 -3.235 ;
        RECT 604.355 -3.565 604.685 -3.235 ;
        RECT 602.995 -3.565 603.325 -3.235 ;
        RECT 601.635 -3.565 601.965 -3.235 ;
        RECT 600.275 -3.565 600.605 -3.235 ;
        RECT 598.915 -3.565 599.245 -3.235 ;
        RECT 597.555 -3.565 597.885 -3.235 ;
        RECT 596.195 -3.565 596.525 -3.235 ;
        RECT 594.835 -3.565 595.165 -3.235 ;
        RECT 593.475 -3.565 593.805 -3.235 ;
        RECT 592.115 -3.565 592.445 -3.235 ;
        RECT 590.755 -3.565 591.085 -3.235 ;
        RECT 589.395 -3.565 589.725 -3.235 ;
        RECT 588.035 -3.565 588.365 -3.235 ;
        RECT 586.675 -3.565 587.005 -3.235 ;
        RECT 585.315 -3.565 585.645 -3.235 ;
        RECT 583.955 -3.565 584.285 -3.235 ;
        RECT 582.595 -3.565 582.925 -3.235 ;
        RECT 581.235 -3.565 581.565 -3.235 ;
        RECT 579.875 -3.565 580.205 -3.235 ;
        RECT 578.515 -3.565 578.845 -3.235 ;
        RECT 577.155 -3.565 577.485 -3.235 ;
        RECT 575.795 -3.565 576.125 -3.235 ;
        RECT 574.435 -3.565 574.765 -3.235 ;
        RECT 573.075 -3.565 573.405 -3.235 ;
        RECT 571.715 -3.565 572.045 -3.235 ;
        RECT 570.355 -3.565 570.685 -3.235 ;
        RECT 568.995 -3.565 569.325 -3.235 ;
        RECT 567.635 -3.565 567.965 -3.235 ;
        RECT 566.275 -3.565 566.605 -3.235 ;
        RECT 564.915 -3.565 565.245 -3.235 ;
        RECT 563.555 -3.565 563.885 -3.235 ;
        RECT 562.195 -3.565 562.525 -3.235 ;
        RECT 560.835 -3.565 561.165 -3.235 ;
        RECT 559.475 -3.565 559.805 -3.235 ;
        RECT 558.115 -3.565 558.445 -3.235 ;
        RECT 556.755 -3.565 557.085 -3.235 ;
        RECT 555.395 -3.565 555.725 -3.235 ;
        RECT 554.035 -3.565 554.365 -3.235 ;
        RECT 552.675 -3.565 553.005 -3.235 ;
        RECT 551.315 -3.565 551.645 -3.235 ;
        RECT 549.955 -3.565 550.285 -3.235 ;
        RECT 548.595 -3.565 548.925 -3.235 ;
        RECT 547.235 -3.565 547.565 -3.235 ;
        RECT 545.875 -3.565 546.205 -3.235 ;
        RECT 544.515 -3.565 544.845 -3.235 ;
        RECT 543.155 -3.565 543.485 -3.235 ;
        RECT 541.795 -3.565 542.125 -3.235 ;
        RECT 540.435 -3.565 540.765 -3.235 ;
        RECT 539.075 -3.565 539.405 -3.235 ;
        RECT 537.715 -3.565 538.045 -3.235 ;
        RECT 536.355 -3.565 536.685 -3.235 ;
        RECT 534.995 -3.565 535.325 -3.235 ;
        RECT 533.635 -3.565 533.965 -3.235 ;
        RECT 532.275 -3.565 532.605 -3.235 ;
        RECT 530.915 -3.565 531.245 -3.235 ;
        RECT 529.555 -3.565 529.885 -3.235 ;
        RECT 528.195 -3.565 528.525 -3.235 ;
        RECT 526.835 -3.565 527.165 -3.235 ;
        RECT 525.475 -3.565 525.805 -3.235 ;
        RECT 524.115 -3.565 524.445 -3.235 ;
        RECT 522.755 -3.565 523.085 -3.235 ;
        RECT 521.395 -3.565 521.725 -3.235 ;
        RECT 520.035 -3.565 520.365 -3.235 ;
        RECT 518.675 -3.565 519.005 -3.235 ;
        RECT 517.315 -3.565 517.645 -3.235 ;
        RECT 515.955 -3.565 516.285 -3.235 ;
        RECT 514.595 -3.565 514.925 -3.235 ;
        RECT 513.235 -3.565 513.565 -3.235 ;
        RECT 511.875 -3.565 512.205 -3.235 ;
        RECT 510.515 -3.565 510.845 -3.235 ;
        RECT 509.155 -3.565 509.485 -3.235 ;
        RECT 507.795 -3.565 508.125 -3.235 ;
        RECT 506.435 -3.565 506.765 -3.235 ;
        RECT 505.075 -3.565 505.405 -3.235 ;
        RECT 503.715 -3.565 504.045 -3.235 ;
        RECT 502.355 -3.565 502.685 -3.235 ;
        RECT 500.995 -3.565 501.325 -3.235 ;
        RECT 499.635 -3.565 499.965 -3.235 ;
        RECT 498.275 -3.565 498.605 -3.235 ;
        RECT 496.915 -3.565 497.245 -3.235 ;
        RECT 495.555 -3.565 495.885 -3.235 ;
        RECT 494.195 -3.565 494.525 -3.235 ;
        RECT 492.835 -3.565 493.165 -3.235 ;
        RECT 491.475 -3.565 491.805 -3.235 ;
        RECT 490.115 -3.565 490.445 -3.235 ;
        RECT 488.755 -3.565 489.085 -3.235 ;
        RECT 487.395 -3.565 487.725 -3.235 ;
        RECT 486.035 -3.565 486.365 -3.235 ;
        RECT 484.675 -3.565 485.005 -3.235 ;
        RECT 483.315 -3.565 483.645 -3.235 ;
        RECT 481.955 -3.565 482.285 -3.235 ;
        RECT 480.595 -3.565 480.925 -3.235 ;
        RECT 479.235 -3.565 479.565 -3.235 ;
        RECT 477.875 -3.565 478.205 -3.235 ;
        RECT 476.515 -3.565 476.845 -3.235 ;
        RECT 475.155 -3.565 475.485 -3.235 ;
        RECT 473.795 -3.565 474.125 -3.235 ;
        RECT 472.435 -3.565 472.765 -3.235 ;
        RECT 471.075 -3.565 471.405 -3.235 ;
        RECT 469.715 -3.565 470.045 -3.235 ;
        RECT 468.355 -3.565 468.685 -3.235 ;
        RECT 466.995 -3.565 467.325 -3.235 ;
        RECT 465.635 -3.565 465.965 -3.235 ;
        RECT 464.275 -3.565 464.605 -3.235 ;
        RECT 462.915 -3.565 463.245 -3.235 ;
        RECT 461.555 -3.565 461.885 -3.235 ;
        RECT 460.195 -3.565 460.525 -3.235 ;
        RECT 458.835 -3.565 459.165 -3.235 ;
        RECT 457.475 -3.565 457.805 -3.235 ;
        RECT 456.115 -3.565 456.445 -3.235 ;
        RECT 454.755 -3.565 455.085 -3.235 ;
        RECT 453.395 -3.565 453.725 -3.235 ;
        RECT 452.035 -3.565 452.365 -3.235 ;
        RECT 450.675 -3.565 451.005 -3.235 ;
        RECT 449.315 -3.565 449.645 -3.235 ;
        RECT 447.955 -3.565 448.285 -3.235 ;
        RECT 446.595 -3.565 446.925 -3.235 ;
        RECT 445.235 -3.565 445.565 -3.235 ;
        RECT 443.875 -3.565 444.205 -3.235 ;
        RECT 442.515 -3.565 442.845 -3.235 ;
        RECT 441.155 -3.565 441.485 -3.235 ;
        RECT 439.795 -3.565 440.125 -3.235 ;
        RECT 438.435 -3.565 438.765 -3.235 ;
        RECT 437.075 -3.565 437.405 -3.235 ;
        RECT 435.715 -3.565 436.045 -3.235 ;
        RECT 434.355 -3.565 434.685 -3.235 ;
        RECT 432.995 -3.565 433.325 -3.235 ;
        RECT 431.635 -3.565 431.965 -3.235 ;
        RECT 430.275 -3.565 430.605 -3.235 ;
        RECT 428.915 -3.565 429.245 -3.235 ;
        RECT 427.555 -3.565 427.885 -3.235 ;
        RECT 426.195 -3.565 426.525 -3.235 ;
        RECT 424.835 -3.565 425.165 -3.235 ;
        RECT 423.475 -3.565 423.805 -3.235 ;
        RECT 422.115 -3.565 422.445 -3.235 ;
        RECT 420.755 -3.565 421.085 -3.235 ;
        RECT 419.395 -3.565 419.725 -3.235 ;
        RECT 418.035 -3.565 418.365 -3.235 ;
        RECT 416.675 -3.565 417.005 -3.235 ;
        RECT 415.315 -3.565 415.645 -3.235 ;
        RECT 413.955 -3.565 414.285 -3.235 ;
        RECT 412.595 -3.565 412.925 -3.235 ;
        RECT 411.235 -3.565 411.565 -3.235 ;
        RECT 409.875 -3.565 410.205 -3.235 ;
        RECT 408.515 -3.565 408.845 -3.235 ;
        RECT 407.155 -3.565 407.485 -3.235 ;
        RECT 405.795 -3.565 406.125 -3.235 ;
        RECT 404.435 -3.565 404.765 -3.235 ;
        RECT 403.075 -3.565 403.405 -3.235 ;
        RECT 401.715 -3.565 402.045 -3.235 ;
        RECT 400.355 -3.565 400.685 -3.235 ;
        RECT 398.995 -3.565 399.325 -3.235 ;
        RECT 397.635 -3.565 397.965 -3.235 ;
        RECT 396.275 -3.565 396.605 -3.235 ;
        RECT 394.915 -3.565 395.245 -3.235 ;
        RECT 393.555 -3.565 393.885 -3.235 ;
        RECT 392.195 -3.565 392.525 -3.235 ;
        RECT 390.835 -3.565 391.165 -3.235 ;
        RECT 389.475 -3.565 389.805 -3.235 ;
        RECT 388.115 -3.565 388.445 -3.235 ;
        RECT 386.755 -3.565 387.085 -3.235 ;
        RECT 385.395 -3.565 385.725 -3.235 ;
        RECT 384.035 -3.565 384.365 -3.235 ;
        RECT 382.675 -3.565 383.005 -3.235 ;
        RECT 381.315 -3.565 381.645 -3.235 ;
        RECT 379.955 -3.565 380.285 -3.235 ;
        RECT 378.595 -3.565 378.925 -3.235 ;
        RECT 377.235 -3.565 377.565 -3.235 ;
        RECT 375.875 -3.565 376.205 -3.235 ;
        RECT 374.515 -3.565 374.845 -3.235 ;
        RECT 373.155 -3.565 373.485 -3.235 ;
        RECT 371.795 -3.565 372.125 -3.235 ;
        RECT 370.435 -3.565 370.765 -3.235 ;
        RECT 369.075 -3.565 369.405 -3.235 ;
        RECT 367.715 -3.565 368.045 -3.235 ;
        RECT 366.355 -3.565 366.685 -3.235 ;
        RECT 364.995 -3.565 365.325 -3.235 ;
        RECT 363.635 -3.565 363.965 -3.235 ;
        RECT 362.275 -3.565 362.605 -3.235 ;
        RECT 360.915 -3.565 361.245 -3.235 ;
        RECT 359.555 -3.565 359.885 -3.235 ;
        RECT 358.195 -3.565 358.525 -3.235 ;
        RECT 356.835 -3.565 357.165 -3.235 ;
        RECT 355.475 -3.565 355.805 -3.235 ;
        RECT 354.115 -3.565 354.445 -3.235 ;
        RECT 352.755 -3.565 353.085 -3.235 ;
        RECT 351.395 -3.565 351.725 -3.235 ;
        RECT 350.035 -3.565 350.365 -3.235 ;
        RECT 348.675 -3.565 349.005 -3.235 ;
        RECT 347.315 -3.565 347.645 -3.235 ;
        RECT 345.955 -3.565 346.285 -3.235 ;
        RECT 344.595 -3.565 344.925 -3.235 ;
        RECT 343.235 -3.565 343.565 -3.235 ;
        RECT 341.875 -3.565 342.205 -3.235 ;
        RECT 340.515 -3.565 340.845 -3.235 ;
        RECT 339.155 -3.565 339.485 -3.235 ;
        RECT 337.795 -3.565 338.125 -3.235 ;
        RECT 336.435 -3.565 336.765 -3.235 ;
        RECT 335.075 -3.565 335.405 -3.235 ;
        RECT 333.715 -3.565 334.045 -3.235 ;
        RECT 332.355 -3.565 332.685 -3.235 ;
        RECT 330.995 -3.565 331.325 -3.235 ;
        RECT 329.635 -3.565 329.965 -3.235 ;
        RECT 328.275 -3.565 328.605 -3.235 ;
        RECT 326.915 -3.565 327.245 -3.235 ;
        RECT 325.555 -3.565 325.885 -3.235 ;
        RECT 324.195 -3.565 324.525 -3.235 ;
        RECT 322.835 -3.565 323.165 -3.235 ;
        RECT 321.475 -3.565 321.805 -3.235 ;
        RECT 320.115 -3.565 320.445 -3.235 ;
        RECT 318.755 -3.565 319.085 -3.235 ;
        RECT 317.395 -3.565 317.725 -3.235 ;
        RECT 316.035 -3.565 316.365 -3.235 ;
        RECT 314.675 -3.565 315.005 -3.235 ;
        RECT 313.315 -3.565 313.645 -3.235 ;
        RECT 311.955 -3.565 312.285 -3.235 ;
        RECT 310.595 -3.565 310.925 -3.235 ;
        RECT 309.235 -3.565 309.565 -3.235 ;
        RECT 307.875 -3.565 308.205 -3.235 ;
        RECT 306.515 -3.565 306.845 -3.235 ;
        RECT 305.155 -3.565 305.485 -3.235 ;
        RECT 303.795 -3.565 304.125 -3.235 ;
        RECT 302.435 -3.565 302.765 -3.235 ;
        RECT 301.075 -3.565 301.405 -3.235 ;
        RECT 299.715 -3.565 300.045 -3.235 ;
        RECT 298.355 -3.565 298.685 -3.235 ;
        RECT 296.995 -3.565 297.325 -3.235 ;
        RECT 295.635 -3.565 295.965 -3.235 ;
        RECT 294.275 -3.565 294.605 -3.235 ;
        RECT 292.915 -3.565 293.245 -3.235 ;
        RECT 291.555 -3.565 291.885 -3.235 ;
        RECT 290.195 -3.565 290.525 -3.235 ;
        RECT 288.835 -3.565 289.165 -3.235 ;
        RECT 287.475 -3.565 287.805 -3.235 ;
        RECT 286.115 -3.565 286.445 -3.235 ;
        RECT 284.755 -3.565 285.085 -3.235 ;
        RECT 283.395 -3.565 283.725 -3.235 ;
        RECT 282.035 -3.565 282.365 -3.235 ;
        RECT 280.675 -3.565 281.005 -3.235 ;
        RECT 279.315 -3.565 279.645 -3.235 ;
        RECT 277.955 -3.565 278.285 -3.235 ;
        RECT 276.595 -3.565 276.925 -3.235 ;
        RECT 275.235 -3.565 275.565 -3.235 ;
        RECT 273.875 -3.565 274.205 -3.235 ;
        RECT 272.515 -3.565 272.845 -3.235 ;
        RECT 271.155 -3.565 271.485 -3.235 ;
        RECT 269.795 -3.565 270.125 -3.235 ;
        RECT 268.435 -3.565 268.765 -3.235 ;
        RECT 267.075 -3.565 267.405 -3.235 ;
        RECT 265.715 -3.565 266.045 -3.235 ;
        RECT 264.355 -3.565 264.685 -3.235 ;
        RECT 262.995 -3.565 263.325 -3.235 ;
        RECT 261.635 -3.565 261.965 -3.235 ;
        RECT 260.275 -3.565 260.605 -3.235 ;
        RECT 258.915 -3.565 259.245 -3.235 ;
        RECT 257.555 -3.565 257.885 -3.235 ;
        RECT 256.195 -3.565 256.525 -3.235 ;
        RECT 254.835 -3.565 255.165 -3.235 ;
        RECT 253.475 -3.565 253.805 -3.235 ;
        RECT 252.115 -3.565 252.445 -3.235 ;
        RECT 250.755 -3.565 251.085 -3.235 ;
        RECT 249.395 -3.565 249.725 -3.235 ;
        RECT 248.035 -3.565 248.365 -3.235 ;
        RECT 246.675 -3.565 247.005 -3.235 ;
        RECT 245.315 -3.565 245.645 -3.235 ;
        RECT 243.955 -3.565 244.285 -3.235 ;
        RECT 242.595 -3.565 242.925 -3.235 ;
        RECT 241.235 -3.565 241.565 -3.235 ;
        RECT 239.875 -3.565 240.205 -3.235 ;
        RECT 238.515 -3.565 238.845 -3.235 ;
        RECT 237.155 -3.565 237.485 -3.235 ;
        RECT 235.795 -3.565 236.125 -3.235 ;
        RECT 234.435 -3.565 234.765 -3.235 ;
        RECT 233.075 -3.565 233.405 -3.235 ;
        RECT 231.715 -3.565 232.045 -3.235 ;
        RECT 230.355 -3.565 230.685 -3.235 ;
        RECT 228.995 -3.565 229.325 -3.235 ;
        RECT 227.635 -3.565 227.965 -3.235 ;
        RECT 226.275 -3.565 226.605 -3.235 ;
        RECT 224.915 -3.565 225.245 -3.235 ;
        RECT 223.555 -3.565 223.885 -3.235 ;
        RECT 222.195 -3.565 222.525 -3.235 ;
        RECT 220.835 -3.565 221.165 -3.235 ;
        RECT 219.475 -3.565 219.805 -3.235 ;
        RECT 218.115 -3.565 218.445 -3.235 ;
        RECT 216.755 -3.565 217.085 -3.235 ;
        RECT 215.395 -3.565 215.725 -3.235 ;
        RECT 214.035 -3.565 214.365 -3.235 ;
        RECT 212.675 -3.565 213.005 -3.235 ;
        RECT 211.315 -3.565 211.645 -3.235 ;
        RECT 209.955 -3.565 210.285 -3.235 ;
        RECT 208.595 -3.565 208.925 -3.235 ;
        RECT 207.235 -3.565 207.565 -3.235 ;
        RECT 205.875 -3.565 206.205 -3.235 ;
        RECT 204.515 -3.565 204.845 -3.235 ;
        RECT 203.155 -3.565 203.485 -3.235 ;
        RECT 201.795 -3.565 202.125 -3.235 ;
        RECT 200.435 -3.565 200.765 -3.235 ;
        RECT 199.075 -3.565 199.405 -3.235 ;
        RECT 197.715 -3.565 198.045 -3.235 ;
        RECT 196.355 -3.565 196.685 -3.235 ;
        RECT 194.995 -3.565 195.325 -3.235 ;
        RECT 193.635 -3.565 193.965 -3.235 ;
        RECT 192.275 -3.565 192.605 -3.235 ;
        RECT 190.915 -3.565 191.245 -3.235 ;
        RECT 189.555 -3.565 189.885 -3.235 ;
        RECT 188.195 -3.565 188.525 -3.235 ;
        RECT 186.835 -3.565 187.165 -3.235 ;
        RECT 185.475 -3.565 185.805 -3.235 ;
        RECT 184.115 -3.565 184.445 -3.235 ;
        RECT 182.755 -3.565 183.085 -3.235 ;
        RECT 181.395 -3.565 181.725 -3.235 ;
        RECT 180.035 -3.565 180.365 -3.235 ;
        RECT 178.675 -3.565 179.005 -3.235 ;
        RECT 177.315 -3.565 177.645 -3.235 ;
        RECT 175.955 -3.565 176.285 -3.235 ;
        RECT 174.595 -3.565 174.925 -3.235 ;
        RECT 173.235 -3.565 173.565 -3.235 ;
        RECT 171.875 -3.565 172.205 -3.235 ;
        RECT 170.515 -3.565 170.845 -3.235 ;
        RECT 169.155 -3.565 169.485 -3.235 ;
        RECT 167.795 -3.565 168.125 -3.235 ;
        RECT 166.435 -3.565 166.765 -3.235 ;
        RECT 165.075 -3.565 165.405 -3.235 ;
        RECT 163.715 -3.565 164.045 -3.235 ;
        RECT 162.355 -3.565 162.685 -3.235 ;
        RECT 160.995 -3.565 161.325 -3.235 ;
        RECT 159.635 -3.565 159.965 -3.235 ;
        RECT 158.275 -3.565 158.605 -3.235 ;
        RECT 156.915 -3.565 157.245 -3.235 ;
        RECT 155.555 -3.565 155.885 -3.235 ;
        RECT 154.195 -3.565 154.525 -3.235 ;
        RECT 152.835 -3.565 153.165 -3.235 ;
        RECT 151.475 -3.565 151.805 -3.235 ;
        RECT 150.115 -3.565 150.445 -3.235 ;
        RECT 148.755 -3.565 149.085 -3.235 ;
        RECT 147.395 -3.565 147.725 -3.235 ;
        RECT 146.035 -3.565 146.365 -3.235 ;
        RECT 144.675 -3.565 145.005 -3.235 ;
        RECT 143.315 -3.565 143.645 -3.235 ;
        RECT 141.955 -3.565 142.285 -3.235 ;
        RECT 140.595 -3.565 140.925 -3.235 ;
        RECT 139.235 -3.565 139.565 -3.235 ;
        RECT 137.875 -3.565 138.205 -3.235 ;
        RECT 678.125 -3.56 954.88 -3.24 ;
        RECT 953.875 -3.565 954.205 -3.235 ;
        RECT 952.515 -3.565 952.845 -3.235 ;
        RECT 951.155 -3.565 951.485 -3.235 ;
        RECT 949.795 -3.565 950.125 -3.235 ;
        RECT 948.435 -3.565 948.765 -3.235 ;
        RECT 947.075 -3.565 947.405 -3.235 ;
        RECT 945.715 -3.565 946.045 -3.235 ;
        RECT 944.355 -3.565 944.685 -3.235 ;
        RECT 942.995 -3.565 943.325 -3.235 ;
        RECT 941.635 -3.565 941.965 -3.235 ;
        RECT 940.275 -3.565 940.605 -3.235 ;
        RECT 938.915 -3.565 939.245 -3.235 ;
        RECT 937.555 -3.565 937.885 -3.235 ;
        RECT 936.195 -3.565 936.525 -3.235 ;
        RECT 934.835 -3.565 935.165 -3.235 ;
        RECT 933.475 -3.565 933.805 -3.235 ;
        RECT 932.115 -3.565 932.445 -3.235 ;
        RECT 930.755 -3.565 931.085 -3.235 ;
        RECT 929.395 -3.565 929.725 -3.235 ;
        RECT 928.035 -3.565 928.365 -3.235 ;
        RECT 926.675 -3.565 927.005 -3.235 ;
        RECT 925.315 -3.565 925.645 -3.235 ;
        RECT 923.955 -3.565 924.285 -3.235 ;
        RECT 922.595 -3.565 922.925 -3.235 ;
        RECT 921.235 -3.565 921.565 -3.235 ;
        RECT 919.875 -3.565 920.205 -3.235 ;
        RECT 918.515 -3.565 918.845 -3.235 ;
        RECT 917.155 -3.565 917.485 -3.235 ;
        RECT 915.795 -3.565 916.125 -3.235 ;
        RECT 914.435 -3.565 914.765 -3.235 ;
        RECT 913.075 -3.565 913.405 -3.235 ;
        RECT 911.715 -3.565 912.045 -3.235 ;
        RECT 910.355 -3.565 910.685 -3.235 ;
        RECT 908.995 -3.565 909.325 -3.235 ;
        RECT 907.635 -3.565 907.965 -3.235 ;
        RECT 906.275 -3.565 906.605 -3.235 ;
        RECT 904.915 -3.565 905.245 -3.235 ;
        RECT 903.555 -3.565 903.885 -3.235 ;
        RECT 902.195 -3.565 902.525 -3.235 ;
        RECT 900.835 -3.565 901.165 -3.235 ;
        RECT 899.475 -3.565 899.805 -3.235 ;
        RECT 898.115 -3.565 898.445 -3.235 ;
        RECT 896.755 -3.565 897.085 -3.235 ;
        RECT 895.395 -3.565 895.725 -3.235 ;
        RECT 894.035 -3.565 894.365 -3.235 ;
        RECT 892.675 -3.565 893.005 -3.235 ;
        RECT 891.315 -3.565 891.645 -3.235 ;
        RECT 889.955 -3.565 890.285 -3.235 ;
        RECT 888.595 -3.565 888.925 -3.235 ;
        RECT 887.235 -3.565 887.565 -3.235 ;
        RECT 885.875 -3.565 886.205 -3.235 ;
        RECT 884.515 -3.565 884.845 -3.235 ;
        RECT 883.155 -3.565 883.485 -3.235 ;
        RECT 881.795 -3.565 882.125 -3.235 ;
        RECT 880.435 -3.565 880.765 -3.235 ;
        RECT 879.075 -3.565 879.405 -3.235 ;
        RECT 877.715 -3.565 878.045 -3.235 ;
        RECT 876.355 -3.565 876.685 -3.235 ;
        RECT 874.995 -3.565 875.325 -3.235 ;
        RECT 873.635 -3.565 873.965 -3.235 ;
        RECT 872.275 -3.565 872.605 -3.235 ;
        RECT 870.915 -3.565 871.245 -3.235 ;
        RECT 869.555 -3.565 869.885 -3.235 ;
        RECT 868.195 -3.565 868.525 -3.235 ;
        RECT 866.835 -3.565 867.165 -3.235 ;
        RECT 865.475 -3.565 865.805 -3.235 ;
        RECT 864.115 -3.565 864.445 -3.235 ;
        RECT 862.755 -3.565 863.085 -3.235 ;
        RECT 861.395 -3.565 861.725 -3.235 ;
        RECT 860.035 -3.565 860.365 -3.235 ;
        RECT 858.675 -3.565 859.005 -3.235 ;
        RECT 857.315 -3.565 857.645 -3.235 ;
        RECT 855.955 -3.565 856.285 -3.235 ;
        RECT 854.595 -3.565 854.925 -3.235 ;
        RECT 853.235 -3.565 853.565 -3.235 ;
        RECT 851.875 -3.565 852.205 -3.235 ;
        RECT 850.515 -3.565 850.845 -3.235 ;
        RECT 849.155 -3.565 849.485 -3.235 ;
        RECT 847.795 -3.565 848.125 -3.235 ;
        RECT 846.435 -3.565 846.765 -3.235 ;
        RECT 845.075 -3.565 845.405 -3.235 ;
        RECT 843.715 -3.565 844.045 -3.235 ;
        RECT 842.355 -3.565 842.685 -3.235 ;
        RECT 840.995 -3.565 841.325 -3.235 ;
        RECT 839.635 -3.565 839.965 -3.235 ;
        RECT 838.275 -3.565 838.605 -3.235 ;
        RECT 836.915 -3.565 837.245 -3.235 ;
        RECT 835.555 -3.565 835.885 -3.235 ;
        RECT 834.195 -3.565 834.525 -3.235 ;
        RECT 832.835 -3.565 833.165 -3.235 ;
        RECT 831.475 -3.565 831.805 -3.235 ;
        RECT 830.115 -3.565 830.445 -3.235 ;
        RECT 828.755 -3.565 829.085 -3.235 ;
        RECT 827.395 -3.565 827.725 -3.235 ;
        RECT 826.035 -3.565 826.365 -3.235 ;
        RECT 824.675 -3.565 825.005 -3.235 ;
        RECT 823.315 -3.565 823.645 -3.235 ;
        RECT 821.955 -3.565 822.285 -3.235 ;
        RECT 820.595 -3.565 820.925 -3.235 ;
        RECT 819.235 -3.565 819.565 -3.235 ;
        RECT 817.875 -3.565 818.205 -3.235 ;
        RECT 816.515 -3.565 816.845 -3.235 ;
        RECT 815.155 -3.565 815.485 -3.235 ;
        RECT 813.795 -3.565 814.125 -3.235 ;
        RECT 812.435 -3.565 812.765 -3.235 ;
        RECT 811.075 -3.565 811.405 -3.235 ;
        RECT 809.715 -3.565 810.045 -3.235 ;
        RECT 808.355 -3.565 808.685 -3.235 ;
        RECT 806.995 -3.565 807.325 -3.235 ;
        RECT 805.635 -3.565 805.965 -3.235 ;
        RECT 804.275 -3.565 804.605 -3.235 ;
        RECT 802.915 -3.565 803.245 -3.235 ;
        RECT 801.555 -3.565 801.885 -3.235 ;
        RECT 800.195 -3.565 800.525 -3.235 ;
        RECT 798.835 -3.565 799.165 -3.235 ;
        RECT 797.475 -3.565 797.805 -3.235 ;
        RECT 796.115 -3.565 796.445 -3.235 ;
        RECT 794.755 -3.565 795.085 -3.235 ;
        RECT 793.395 -3.565 793.725 -3.235 ;
        RECT 792.035 -3.565 792.365 -3.235 ;
        RECT 790.675 -3.565 791.005 -3.235 ;
        RECT 789.315 -3.565 789.645 -3.235 ;
        RECT 787.955 -3.565 788.285 -3.235 ;
        RECT 786.595 -3.565 786.925 -3.235 ;
        RECT 785.235 -3.565 785.565 -3.235 ;
        RECT 783.875 -3.565 784.205 -3.235 ;
        RECT 782.515 -3.565 782.845 -3.235 ;
        RECT 781.155 -3.565 781.485 -3.235 ;
        RECT 779.795 -3.565 780.125 -3.235 ;
        RECT 778.435 -3.565 778.765 -3.235 ;
        RECT 777.075 -3.565 777.405 -3.235 ;
        RECT 775.715 -3.565 776.045 -3.235 ;
        RECT 774.355 -3.565 774.685 -3.235 ;
        RECT 772.995 -3.565 773.325 -3.235 ;
        RECT 771.635 -3.565 771.965 -3.235 ;
        RECT 770.275 -3.565 770.605 -3.235 ;
        RECT 768.915 -3.565 769.245 -3.235 ;
        RECT 767.555 -3.565 767.885 -3.235 ;
        RECT 766.195 -3.565 766.525 -3.235 ;
        RECT 764.835 -3.565 765.165 -3.235 ;
        RECT 763.475 -3.565 763.805 -3.235 ;
        RECT 762.115 -3.565 762.445 -3.235 ;
        RECT 760.755 -3.565 761.085 -3.235 ;
        RECT 759.395 -3.565 759.725 -3.235 ;
        RECT 758.035 -3.565 758.365 -3.235 ;
        RECT 756.675 -3.565 757.005 -3.235 ;
        RECT 755.315 -3.565 755.645 -3.235 ;
        RECT 753.955 -3.565 754.285 -3.235 ;
        RECT 752.595 -3.565 752.925 -3.235 ;
        RECT 751.235 -3.565 751.565 -3.235 ;
        RECT 749.875 -3.565 750.205 -3.235 ;
        RECT 748.515 -3.565 748.845 -3.235 ;
        RECT 747.155 -3.565 747.485 -3.235 ;
        RECT 745.795 -3.565 746.125 -3.235 ;
        RECT 744.435 -3.565 744.765 -3.235 ;
        RECT 743.075 -3.565 743.405 -3.235 ;
        RECT 741.715 -3.565 742.045 -3.235 ;
        RECT 740.355 -3.565 740.685 -3.235 ;
        RECT 738.995 -3.565 739.325 -3.235 ;
        RECT 737.635 -3.565 737.965 -3.235 ;
        RECT 736.275 -3.565 736.605 -3.235 ;
        RECT 734.915 -3.565 735.245 -3.235 ;
        RECT 733.555 -3.565 733.885 -3.235 ;
        RECT 732.195 -3.565 732.525 -3.235 ;
        RECT 730.835 -3.565 731.165 -3.235 ;
        RECT 729.475 -3.565 729.805 -3.235 ;
        RECT 728.115 -3.565 728.445 -3.235 ;
        RECT 726.755 -3.565 727.085 -3.235 ;
        RECT 725.395 -3.565 725.725 -3.235 ;
        RECT 724.035 -3.565 724.365 -3.235 ;
        RECT 722.675 -3.565 723.005 -3.235 ;
        RECT 721.315 -3.565 721.645 -3.235 ;
        RECT 719.955 -3.565 720.285 -3.235 ;
        RECT 718.595 -3.565 718.925 -3.235 ;
        RECT 717.235 -3.565 717.565 -3.235 ;
        RECT 715.875 -3.565 716.205 -3.235 ;
        RECT 714.515 -3.565 714.845 -3.235 ;
        RECT 713.155 -3.565 713.485 -3.235 ;
        RECT 711.795 -3.565 712.125 -3.235 ;
        RECT 710.435 -3.565 710.765 -3.235 ;
        RECT 709.075 -3.565 709.405 -3.235 ;
        RECT 707.715 -3.565 708.045 -3.235 ;
        RECT 706.355 -3.565 706.685 -3.235 ;
        RECT 704.995 -3.565 705.325 -3.235 ;
        RECT 703.635 -3.565 703.965 -3.235 ;
        RECT 702.275 -3.565 702.605 -3.235 ;
        RECT 700.915 -3.565 701.245 -3.235 ;
        RECT 699.555 -3.565 699.885 -3.235 ;
        RECT 698.195 -3.565 698.525 -3.235 ;
        RECT 696.835 -3.565 697.165 -3.235 ;
        RECT 695.475 -3.565 695.805 -3.235 ;
        RECT 694.115 -3.565 694.445 -3.235 ;
        RECT 692.755 -3.565 693.085 -3.235 ;
        RECT 691.395 -3.565 691.725 -3.235 ;
        RECT 690.035 -3.565 690.365 -3.235 ;
        RECT 688.675 -3.565 689.005 -3.235 ;
        RECT 687.315 -3.565 687.645 -3.235 ;
        RECT 685.955 -3.565 686.285 -3.235 ;
        RECT 684.595 -3.565 684.925 -3.235 ;
        RECT 683.235 -3.565 683.565 -3.235 ;
        RECT 681.875 -3.565 682.205 -3.235 ;
        RECT 680.515 -3.565 680.845 -3.235 ;
        RECT 679.155 -3.565 679.485 -3.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.795 0.515 678.125 0.845 ;
        RECT -1.52 0.52 678.125 0.84 ;
        RECT 676.435 0.515 676.765 0.845 ;
        RECT 675.075 0.515 675.405 0.845 ;
        RECT 673.715 0.515 674.045 0.845 ;
        RECT 672.355 0.515 672.685 0.845 ;
        RECT 670.995 0.515 671.325 0.845 ;
        RECT 669.635 0.515 669.965 0.845 ;
        RECT 668.275 0.515 668.605 0.845 ;
        RECT 666.915 0.515 667.245 0.845 ;
        RECT 665.555 0.515 665.885 0.845 ;
        RECT 664.195 0.515 664.525 0.845 ;
        RECT 662.835 0.515 663.165 0.845 ;
        RECT 661.475 0.515 661.805 0.845 ;
        RECT 660.115 0.515 660.445 0.845 ;
        RECT 658.755 0.515 659.085 0.845 ;
        RECT 657.395 0.515 657.725 0.845 ;
        RECT 656.035 0.515 656.365 0.845 ;
        RECT 654.675 0.515 655.005 0.845 ;
        RECT 653.315 0.515 653.645 0.845 ;
        RECT 651.955 0.515 652.285 0.845 ;
        RECT 650.595 0.515 650.925 0.845 ;
        RECT 649.235 0.515 649.565 0.845 ;
        RECT 647.875 0.515 648.205 0.845 ;
        RECT 646.515 0.515 646.845 0.845 ;
        RECT 645.155 0.515 645.485 0.845 ;
        RECT 643.795 0.515 644.125 0.845 ;
        RECT 642.435 0.515 642.765 0.845 ;
        RECT 641.075 0.515 641.405 0.845 ;
        RECT 639.715 0.515 640.045 0.845 ;
        RECT 638.355 0.515 638.685 0.845 ;
        RECT 636.995 0.515 637.325 0.845 ;
        RECT 635.635 0.515 635.965 0.845 ;
        RECT 634.275 0.515 634.605 0.845 ;
        RECT 632.915 0.515 633.245 0.845 ;
        RECT 631.555 0.515 631.885 0.845 ;
        RECT 630.195 0.515 630.525 0.845 ;
        RECT 628.835 0.515 629.165 0.845 ;
        RECT 627.475 0.515 627.805 0.845 ;
        RECT 626.115 0.515 626.445 0.845 ;
        RECT 624.755 0.515 625.085 0.845 ;
        RECT 623.395 0.515 623.725 0.845 ;
        RECT 622.035 0.515 622.365 0.845 ;
        RECT 620.675 0.515 621.005 0.845 ;
        RECT 619.315 0.515 619.645 0.845 ;
        RECT 617.955 0.515 618.285 0.845 ;
        RECT 616.595 0.515 616.925 0.845 ;
        RECT 615.235 0.515 615.565 0.845 ;
        RECT 613.875 0.515 614.205 0.845 ;
        RECT 612.515 0.515 612.845 0.845 ;
        RECT 611.155 0.515 611.485 0.845 ;
        RECT 609.795 0.515 610.125 0.845 ;
        RECT 608.435 0.515 608.765 0.845 ;
        RECT 607.075 0.515 607.405 0.845 ;
        RECT 605.715 0.515 606.045 0.845 ;
        RECT 604.355 0.515 604.685 0.845 ;
        RECT 602.995 0.515 603.325 0.845 ;
        RECT 601.635 0.515 601.965 0.845 ;
        RECT 600.275 0.515 600.605 0.845 ;
        RECT 598.915 0.515 599.245 0.845 ;
        RECT 597.555 0.515 597.885 0.845 ;
        RECT 596.195 0.515 596.525 0.845 ;
        RECT 594.835 0.515 595.165 0.845 ;
        RECT 593.475 0.515 593.805 0.845 ;
        RECT 592.115 0.515 592.445 0.845 ;
        RECT 590.755 0.515 591.085 0.845 ;
        RECT 589.395 0.515 589.725 0.845 ;
        RECT 588.035 0.515 588.365 0.845 ;
        RECT 586.675 0.515 587.005 0.845 ;
        RECT 585.315 0.515 585.645 0.845 ;
        RECT 583.955 0.515 584.285 0.845 ;
        RECT 582.595 0.515 582.925 0.845 ;
        RECT 581.235 0.515 581.565 0.845 ;
        RECT 579.875 0.515 580.205 0.845 ;
        RECT 578.515 0.515 578.845 0.845 ;
        RECT 577.155 0.515 577.485 0.845 ;
        RECT 575.795 0.515 576.125 0.845 ;
        RECT 574.435 0.515 574.765 0.845 ;
        RECT 573.075 0.515 573.405 0.845 ;
        RECT 571.715 0.515 572.045 0.845 ;
        RECT 570.355 0.515 570.685 0.845 ;
        RECT 568.995 0.515 569.325 0.845 ;
        RECT 567.635 0.515 567.965 0.845 ;
        RECT 566.275 0.515 566.605 0.845 ;
        RECT 564.915 0.515 565.245 0.845 ;
        RECT 563.555 0.515 563.885 0.845 ;
        RECT 562.195 0.515 562.525 0.845 ;
        RECT 560.835 0.515 561.165 0.845 ;
        RECT 559.475 0.515 559.805 0.845 ;
        RECT 558.115 0.515 558.445 0.845 ;
        RECT 556.755 0.515 557.085 0.845 ;
        RECT 555.395 0.515 555.725 0.845 ;
        RECT 554.035 0.515 554.365 0.845 ;
        RECT 552.675 0.515 553.005 0.845 ;
        RECT 551.315 0.515 551.645 0.845 ;
        RECT 549.955 0.515 550.285 0.845 ;
        RECT 548.595 0.515 548.925 0.845 ;
        RECT 547.235 0.515 547.565 0.845 ;
        RECT 545.875 0.515 546.205 0.845 ;
        RECT 544.515 0.515 544.845 0.845 ;
        RECT 543.155 0.515 543.485 0.845 ;
        RECT 541.795 0.515 542.125 0.845 ;
        RECT 540.435 0.515 540.765 0.845 ;
        RECT 539.075 0.515 539.405 0.845 ;
        RECT 537.715 0.515 538.045 0.845 ;
        RECT 536.355 0.515 536.685 0.845 ;
        RECT 534.995 0.515 535.325 0.845 ;
        RECT 533.635 0.515 533.965 0.845 ;
        RECT 532.275 0.515 532.605 0.845 ;
        RECT 530.915 0.515 531.245 0.845 ;
        RECT 529.555 0.515 529.885 0.845 ;
        RECT 528.195 0.515 528.525 0.845 ;
        RECT 526.835 0.515 527.165 0.845 ;
        RECT 525.475 0.515 525.805 0.845 ;
        RECT 524.115 0.515 524.445 0.845 ;
        RECT 522.755 0.515 523.085 0.845 ;
        RECT 521.395 0.515 521.725 0.845 ;
        RECT 520.035 0.515 520.365 0.845 ;
        RECT 518.675 0.515 519.005 0.845 ;
        RECT 517.315 0.515 517.645 0.845 ;
        RECT 515.955 0.515 516.285 0.845 ;
        RECT 514.595 0.515 514.925 0.845 ;
        RECT 513.235 0.515 513.565 0.845 ;
        RECT 511.875 0.515 512.205 0.845 ;
        RECT 510.515 0.515 510.845 0.845 ;
        RECT 509.155 0.515 509.485 0.845 ;
        RECT 507.795 0.515 508.125 0.845 ;
        RECT 506.435 0.515 506.765 0.845 ;
        RECT 505.075 0.515 505.405 0.845 ;
        RECT 503.715 0.515 504.045 0.845 ;
        RECT 502.355 0.515 502.685 0.845 ;
        RECT 500.995 0.515 501.325 0.845 ;
        RECT 499.635 0.515 499.965 0.845 ;
        RECT 498.275 0.515 498.605 0.845 ;
        RECT 496.915 0.515 497.245 0.845 ;
        RECT 495.555 0.515 495.885 0.845 ;
        RECT 494.195 0.515 494.525 0.845 ;
        RECT 492.835 0.515 493.165 0.845 ;
        RECT 491.475 0.515 491.805 0.845 ;
        RECT 490.115 0.515 490.445 0.845 ;
        RECT 488.755 0.515 489.085 0.845 ;
        RECT 487.395 0.515 487.725 0.845 ;
        RECT 486.035 0.515 486.365 0.845 ;
        RECT 484.675 0.515 485.005 0.845 ;
        RECT 483.315 0.515 483.645 0.845 ;
        RECT 481.955 0.515 482.285 0.845 ;
        RECT 480.595 0.515 480.925 0.845 ;
        RECT 479.235 0.515 479.565 0.845 ;
        RECT 477.875 0.515 478.205 0.845 ;
        RECT 476.515 0.515 476.845 0.845 ;
        RECT 475.155 0.515 475.485 0.845 ;
        RECT 473.795 0.515 474.125 0.845 ;
        RECT 472.435 0.515 472.765 0.845 ;
        RECT 471.075 0.515 471.405 0.845 ;
        RECT 469.715 0.515 470.045 0.845 ;
        RECT 468.355 0.515 468.685 0.845 ;
        RECT 466.995 0.515 467.325 0.845 ;
        RECT 465.635 0.515 465.965 0.845 ;
        RECT 464.275 0.515 464.605 0.845 ;
        RECT 462.915 0.515 463.245 0.845 ;
        RECT 461.555 0.515 461.885 0.845 ;
        RECT 460.195 0.515 460.525 0.845 ;
        RECT 458.835 0.515 459.165 0.845 ;
        RECT 457.475 0.515 457.805 0.845 ;
        RECT 456.115 0.515 456.445 0.845 ;
        RECT 454.755 0.515 455.085 0.845 ;
        RECT 453.395 0.515 453.725 0.845 ;
        RECT 452.035 0.515 452.365 0.845 ;
        RECT 450.675 0.515 451.005 0.845 ;
        RECT 449.315 0.515 449.645 0.845 ;
        RECT 447.955 0.515 448.285 0.845 ;
        RECT 446.595 0.515 446.925 0.845 ;
        RECT 445.235 0.515 445.565 0.845 ;
        RECT 443.875 0.515 444.205 0.845 ;
        RECT 442.515 0.515 442.845 0.845 ;
        RECT 441.155 0.515 441.485 0.845 ;
        RECT 439.795 0.515 440.125 0.845 ;
        RECT 438.435 0.515 438.765 0.845 ;
        RECT 437.075 0.515 437.405 0.845 ;
        RECT 435.715 0.515 436.045 0.845 ;
        RECT 434.355 0.515 434.685 0.845 ;
        RECT 432.995 0.515 433.325 0.845 ;
        RECT 431.635 0.515 431.965 0.845 ;
        RECT 430.275 0.515 430.605 0.845 ;
        RECT 428.915 0.515 429.245 0.845 ;
        RECT 427.555 0.515 427.885 0.845 ;
        RECT 426.195 0.515 426.525 0.845 ;
        RECT 424.835 0.515 425.165 0.845 ;
        RECT 423.475 0.515 423.805 0.845 ;
        RECT 422.115 0.515 422.445 0.845 ;
        RECT 420.755 0.515 421.085 0.845 ;
        RECT 419.395 0.515 419.725 0.845 ;
        RECT 418.035 0.515 418.365 0.845 ;
        RECT 416.675 0.515 417.005 0.845 ;
        RECT 415.315 0.515 415.645 0.845 ;
        RECT 413.955 0.515 414.285 0.845 ;
        RECT 412.595 0.515 412.925 0.845 ;
        RECT 411.235 0.515 411.565 0.845 ;
        RECT 409.875 0.515 410.205 0.845 ;
        RECT 408.515 0.515 408.845 0.845 ;
        RECT 407.155 0.515 407.485 0.845 ;
        RECT 405.795 0.515 406.125 0.845 ;
        RECT 404.435 0.515 404.765 0.845 ;
        RECT 403.075 0.515 403.405 0.845 ;
        RECT 401.715 0.515 402.045 0.845 ;
        RECT 400.355 0.515 400.685 0.845 ;
        RECT 398.995 0.515 399.325 0.845 ;
        RECT 397.635 0.515 397.965 0.845 ;
        RECT 396.275 0.515 396.605 0.845 ;
        RECT 394.915 0.515 395.245 0.845 ;
        RECT 393.555 0.515 393.885 0.845 ;
        RECT 392.195 0.515 392.525 0.845 ;
        RECT 390.835 0.515 391.165 0.845 ;
        RECT 389.475 0.515 389.805 0.845 ;
        RECT 388.115 0.515 388.445 0.845 ;
        RECT 386.755 0.515 387.085 0.845 ;
        RECT 385.395 0.515 385.725 0.845 ;
        RECT 384.035 0.515 384.365 0.845 ;
        RECT 382.675 0.515 383.005 0.845 ;
        RECT 381.315 0.515 381.645 0.845 ;
        RECT 379.955 0.515 380.285 0.845 ;
        RECT 378.595 0.515 378.925 0.845 ;
        RECT 377.235 0.515 377.565 0.845 ;
        RECT 375.875 0.515 376.205 0.845 ;
        RECT 374.515 0.515 374.845 0.845 ;
        RECT 373.155 0.515 373.485 0.845 ;
        RECT 371.795 0.515 372.125 0.845 ;
        RECT 370.435 0.515 370.765 0.845 ;
        RECT 369.075 0.515 369.405 0.845 ;
        RECT 367.715 0.515 368.045 0.845 ;
        RECT 366.355 0.515 366.685 0.845 ;
        RECT 364.995 0.515 365.325 0.845 ;
        RECT 363.635 0.515 363.965 0.845 ;
        RECT 362.275 0.515 362.605 0.845 ;
        RECT 360.915 0.515 361.245 0.845 ;
        RECT 359.555 0.515 359.885 0.845 ;
        RECT 358.195 0.515 358.525 0.845 ;
        RECT 356.835 0.515 357.165 0.845 ;
        RECT 355.475 0.515 355.805 0.845 ;
        RECT 354.115 0.515 354.445 0.845 ;
        RECT 352.755 0.515 353.085 0.845 ;
        RECT 351.395 0.515 351.725 0.845 ;
        RECT 350.035 0.515 350.365 0.845 ;
        RECT 348.675 0.515 349.005 0.845 ;
        RECT 347.315 0.515 347.645 0.845 ;
        RECT 345.955 0.515 346.285 0.845 ;
        RECT 344.595 0.515 344.925 0.845 ;
        RECT 343.235 0.515 343.565 0.845 ;
        RECT 341.875 0.515 342.205 0.845 ;
        RECT 340.515 0.515 340.845 0.845 ;
        RECT 339.155 0.515 339.485 0.845 ;
        RECT 337.795 0.515 338.125 0.845 ;
        RECT 336.435 0.515 336.765 0.845 ;
        RECT 335.075 0.515 335.405 0.845 ;
        RECT 333.715 0.515 334.045 0.845 ;
        RECT 332.355 0.515 332.685 0.845 ;
        RECT 330.995 0.515 331.325 0.845 ;
        RECT 329.635 0.515 329.965 0.845 ;
        RECT 328.275 0.515 328.605 0.845 ;
        RECT 326.915 0.515 327.245 0.845 ;
        RECT 325.555 0.515 325.885 0.845 ;
        RECT 324.195 0.515 324.525 0.845 ;
        RECT 322.835 0.515 323.165 0.845 ;
        RECT 321.475 0.515 321.805 0.845 ;
        RECT 320.115 0.515 320.445 0.845 ;
        RECT 318.755 0.515 319.085 0.845 ;
        RECT 317.395 0.515 317.725 0.845 ;
        RECT 316.035 0.515 316.365 0.845 ;
        RECT 314.675 0.515 315.005 0.845 ;
        RECT 313.315 0.515 313.645 0.845 ;
        RECT 311.955 0.515 312.285 0.845 ;
        RECT 310.595 0.515 310.925 0.845 ;
        RECT 309.235 0.515 309.565 0.845 ;
        RECT 307.875 0.515 308.205 0.845 ;
        RECT 306.515 0.515 306.845 0.845 ;
        RECT 305.155 0.515 305.485 0.845 ;
        RECT 303.795 0.515 304.125 0.845 ;
        RECT 302.435 0.515 302.765 0.845 ;
        RECT 301.075 0.515 301.405 0.845 ;
        RECT 299.715 0.515 300.045 0.845 ;
        RECT 298.355 0.515 298.685 0.845 ;
        RECT 296.995 0.515 297.325 0.845 ;
        RECT 295.635 0.515 295.965 0.845 ;
        RECT 294.275 0.515 294.605 0.845 ;
        RECT 292.915 0.515 293.245 0.845 ;
        RECT 291.555 0.515 291.885 0.845 ;
        RECT 290.195 0.515 290.525 0.845 ;
        RECT 288.835 0.515 289.165 0.845 ;
        RECT 287.475 0.515 287.805 0.845 ;
        RECT 286.115 0.515 286.445 0.845 ;
        RECT 284.755 0.515 285.085 0.845 ;
        RECT 283.395 0.515 283.725 0.845 ;
        RECT 282.035 0.515 282.365 0.845 ;
        RECT 280.675 0.515 281.005 0.845 ;
        RECT 279.315 0.515 279.645 0.845 ;
        RECT 277.955 0.515 278.285 0.845 ;
        RECT 276.595 0.515 276.925 0.845 ;
        RECT 275.235 0.515 275.565 0.845 ;
        RECT 273.875 0.515 274.205 0.845 ;
        RECT 272.515 0.515 272.845 0.845 ;
        RECT 271.155 0.515 271.485 0.845 ;
        RECT 269.795 0.515 270.125 0.845 ;
        RECT 268.435 0.515 268.765 0.845 ;
        RECT 267.075 0.515 267.405 0.845 ;
        RECT 265.715 0.515 266.045 0.845 ;
        RECT 264.355 0.515 264.685 0.845 ;
        RECT 262.995 0.515 263.325 0.845 ;
        RECT 261.635 0.515 261.965 0.845 ;
        RECT 260.275 0.515 260.605 0.845 ;
        RECT 258.915 0.515 259.245 0.845 ;
        RECT 257.555 0.515 257.885 0.845 ;
        RECT 256.195 0.515 256.525 0.845 ;
        RECT 254.835 0.515 255.165 0.845 ;
        RECT 253.475 0.515 253.805 0.845 ;
        RECT 252.115 0.515 252.445 0.845 ;
        RECT 250.755 0.515 251.085 0.845 ;
        RECT 249.395 0.515 249.725 0.845 ;
        RECT 248.035 0.515 248.365 0.845 ;
        RECT 246.675 0.515 247.005 0.845 ;
        RECT 245.315 0.515 245.645 0.845 ;
        RECT 243.955 0.515 244.285 0.845 ;
        RECT 242.595 0.515 242.925 0.845 ;
        RECT 241.235 0.515 241.565 0.845 ;
        RECT 239.875 0.515 240.205 0.845 ;
        RECT 238.515 0.515 238.845 0.845 ;
        RECT 237.155 0.515 237.485 0.845 ;
        RECT 235.795 0.515 236.125 0.845 ;
        RECT 234.435 0.515 234.765 0.845 ;
        RECT 233.075 0.515 233.405 0.845 ;
        RECT 231.715 0.515 232.045 0.845 ;
        RECT 230.355 0.515 230.685 0.845 ;
        RECT 228.995 0.515 229.325 0.845 ;
        RECT 227.635 0.515 227.965 0.845 ;
        RECT 226.275 0.515 226.605 0.845 ;
        RECT 224.915 0.515 225.245 0.845 ;
        RECT 223.555 0.515 223.885 0.845 ;
        RECT 222.195 0.515 222.525 0.845 ;
        RECT 220.835 0.515 221.165 0.845 ;
        RECT 219.475 0.515 219.805 0.845 ;
        RECT 218.115 0.515 218.445 0.845 ;
        RECT 216.755 0.515 217.085 0.845 ;
        RECT 215.395 0.515 215.725 0.845 ;
        RECT 214.035 0.515 214.365 0.845 ;
        RECT 212.675 0.515 213.005 0.845 ;
        RECT 211.315 0.515 211.645 0.845 ;
        RECT 209.955 0.515 210.285 0.845 ;
        RECT 208.595 0.515 208.925 0.845 ;
        RECT 207.235 0.515 207.565 0.845 ;
        RECT 205.875 0.515 206.205 0.845 ;
        RECT 204.515 0.515 204.845 0.845 ;
        RECT 203.155 0.515 203.485 0.845 ;
        RECT 201.795 0.515 202.125 0.845 ;
        RECT 200.435 0.515 200.765 0.845 ;
        RECT 199.075 0.515 199.405 0.845 ;
        RECT 197.715 0.515 198.045 0.845 ;
        RECT 196.355 0.515 196.685 0.845 ;
        RECT 194.995 0.515 195.325 0.845 ;
        RECT 193.635 0.515 193.965 0.845 ;
        RECT 192.275 0.515 192.605 0.845 ;
        RECT 190.915 0.515 191.245 0.845 ;
        RECT 189.555 0.515 189.885 0.845 ;
        RECT 188.195 0.515 188.525 0.845 ;
        RECT 186.835 0.515 187.165 0.845 ;
        RECT 185.475 0.515 185.805 0.845 ;
        RECT 184.115 0.515 184.445 0.845 ;
        RECT 182.755 0.515 183.085 0.845 ;
        RECT 181.395 0.515 181.725 0.845 ;
        RECT 180.035 0.515 180.365 0.845 ;
        RECT 178.675 0.515 179.005 0.845 ;
        RECT 177.315 0.515 177.645 0.845 ;
        RECT 175.955 0.515 176.285 0.845 ;
        RECT 174.595 0.515 174.925 0.845 ;
        RECT 173.235 0.515 173.565 0.845 ;
        RECT 171.875 0.515 172.205 0.845 ;
        RECT 170.515 0.515 170.845 0.845 ;
        RECT 169.155 0.515 169.485 0.845 ;
        RECT 167.795 0.515 168.125 0.845 ;
        RECT 166.435 0.515 166.765 0.845 ;
        RECT 165.075 0.515 165.405 0.845 ;
        RECT 163.715 0.515 164.045 0.845 ;
        RECT 162.355 0.515 162.685 0.845 ;
        RECT 160.995 0.515 161.325 0.845 ;
        RECT 159.635 0.515 159.965 0.845 ;
        RECT 158.275 0.515 158.605 0.845 ;
        RECT 156.915 0.515 157.245 0.845 ;
        RECT 155.555 0.515 155.885 0.845 ;
        RECT 154.195 0.515 154.525 0.845 ;
        RECT 152.835 0.515 153.165 0.845 ;
        RECT 151.475 0.515 151.805 0.845 ;
        RECT 150.115 0.515 150.445 0.845 ;
        RECT 148.755 0.515 149.085 0.845 ;
        RECT 147.395 0.515 147.725 0.845 ;
        RECT 146.035 0.515 146.365 0.845 ;
        RECT 144.675 0.515 145.005 0.845 ;
        RECT 143.315 0.515 143.645 0.845 ;
        RECT 141.955 0.515 142.285 0.845 ;
        RECT 140.595 0.515 140.925 0.845 ;
        RECT 139.235 0.515 139.565 0.845 ;
        RECT 137.875 0.515 138.205 0.845 ;
        RECT 136.515 0.515 136.845 0.845 ;
        RECT 135.155 0.515 135.485 0.845 ;
        RECT 133.795 0.515 134.125 0.845 ;
        RECT 132.435 0.515 132.765 0.845 ;
        RECT 131.075 0.515 131.405 0.845 ;
        RECT 129.715 0.515 130.045 0.845 ;
        RECT 128.355 0.515 128.685 0.845 ;
        RECT 126.995 0.515 127.325 0.845 ;
        RECT 125.635 0.515 125.965 0.845 ;
        RECT 124.275 0.515 124.605 0.845 ;
        RECT 122.915 0.515 123.245 0.845 ;
        RECT 121.555 0.515 121.885 0.845 ;
        RECT 120.195 0.515 120.525 0.845 ;
        RECT 118.835 0.515 119.165 0.845 ;
        RECT 117.475 0.515 117.805 0.845 ;
        RECT 116.115 0.515 116.445 0.845 ;
        RECT 114.755 0.515 115.085 0.845 ;
        RECT 113.395 0.515 113.725 0.845 ;
        RECT 112.035 0.515 112.365 0.845 ;
        RECT 110.675 0.515 111.005 0.845 ;
        RECT 109.315 0.515 109.645 0.845 ;
        RECT 107.955 0.515 108.285 0.845 ;
        RECT 106.595 0.515 106.925 0.845 ;
        RECT 105.235 0.515 105.565 0.845 ;
        RECT 103.875 0.515 104.205 0.845 ;
        RECT 102.515 0.515 102.845 0.845 ;
        RECT 101.155 0.515 101.485 0.845 ;
        RECT 99.795 0.515 100.125 0.845 ;
        RECT 98.435 0.515 98.765 0.845 ;
        RECT 97.075 0.515 97.405 0.845 ;
        RECT 95.715 0.515 96.045 0.845 ;
        RECT 94.355 0.515 94.685 0.845 ;
        RECT 92.995 0.515 93.325 0.845 ;
        RECT 91.635 0.515 91.965 0.845 ;
        RECT 90.275 0.515 90.605 0.845 ;
        RECT 88.915 0.515 89.245 0.845 ;
        RECT 87.555 0.515 87.885 0.845 ;
        RECT 86.195 0.515 86.525 0.845 ;
        RECT 84.835 0.515 85.165 0.845 ;
        RECT 83.475 0.515 83.805 0.845 ;
        RECT 82.115 0.515 82.445 0.845 ;
        RECT 80.755 0.515 81.085 0.845 ;
        RECT 79.395 0.515 79.725 0.845 ;
        RECT 78.035 0.515 78.365 0.845 ;
        RECT 76.675 0.515 77.005 0.845 ;
        RECT 75.315 0.515 75.645 0.845 ;
        RECT 73.955 0.515 74.285 0.845 ;
        RECT 72.595 0.515 72.925 0.845 ;
        RECT 71.235 0.515 71.565 0.845 ;
        RECT 69.875 0.515 70.205 0.845 ;
        RECT 68.515 0.515 68.845 0.845 ;
        RECT 67.155 0.515 67.485 0.845 ;
        RECT 65.795 0.515 66.125 0.845 ;
        RECT 64.435 0.515 64.765 0.845 ;
        RECT 63.075 0.515 63.405 0.845 ;
        RECT 61.715 0.515 62.045 0.845 ;
        RECT 60.355 0.515 60.685 0.845 ;
        RECT 58.995 0.515 59.325 0.845 ;
        RECT 57.635 0.515 57.965 0.845 ;
        RECT 56.275 0.515 56.605 0.845 ;
        RECT 54.915 0.515 55.245 0.845 ;
        RECT 53.555 0.515 53.885 0.845 ;
        RECT 52.195 0.515 52.525 0.845 ;
        RECT 50.835 0.515 51.165 0.845 ;
        RECT 49.475 0.515 49.805 0.845 ;
        RECT 48.115 0.515 48.445 0.845 ;
        RECT 46.755 0.515 47.085 0.845 ;
        RECT 45.395 0.515 45.725 0.845 ;
        RECT 44.035 0.515 44.365 0.845 ;
        RECT 42.675 0.515 43.005 0.845 ;
        RECT 41.315 0.515 41.645 0.845 ;
        RECT 39.955 0.515 40.285 0.845 ;
        RECT 38.595 0.515 38.925 0.845 ;
        RECT 37.235 0.515 37.565 0.845 ;
        RECT 35.875 0.515 36.205 0.845 ;
        RECT 34.515 0.515 34.845 0.845 ;
        RECT 33.155 0.515 33.485 0.845 ;
        RECT 31.795 0.515 32.125 0.845 ;
        RECT 30.435 0.515 30.765 0.845 ;
        RECT 29.075 0.515 29.405 0.845 ;
        RECT 27.715 0.515 28.045 0.845 ;
        RECT 26.355 0.515 26.685 0.845 ;
        RECT 24.995 0.515 25.325 0.845 ;
        RECT 23.635 0.515 23.965 0.845 ;
        RECT 22.275 0.515 22.605 0.845 ;
        RECT 20.915 0.515 21.245 0.845 ;
        RECT 19.555 0.515 19.885 0.845 ;
        RECT 18.195 0.515 18.525 0.845 ;
        RECT 16.835 0.515 17.165 0.845 ;
        RECT 15.475 0.515 15.805 0.845 ;
        RECT 14.115 0.515 14.445 0.845 ;
        RECT 12.755 0.515 13.085 0.845 ;
        RECT 11.395 0.515 11.725 0.845 ;
        RECT 10.035 0.515 10.365 0.845 ;
        RECT 8.675 0.515 9.005 0.845 ;
        RECT 7.315 0.515 7.645 0.845 ;
        RECT 5.955 0.515 6.285 0.845 ;
        RECT 4.595 0.515 4.925 0.845 ;
        RECT 3.235 0.515 3.565 0.845 ;
        RECT 1.875 0.515 2.205 0.845 ;
        RECT 0.515 0.515 0.845 0.845 ;
        RECT -0.845 0.515 -0.515 0.845 ;
        RECT 678.125 0.52 954.88 0.84 ;
        RECT 953.875 0.515 954.205 0.845 ;
        RECT 952.515 0.515 952.845 0.845 ;
        RECT 951.155 0.515 951.485 0.845 ;
        RECT 949.795 0.515 950.125 0.845 ;
        RECT 948.435 0.515 948.765 0.845 ;
        RECT 947.075 0.515 947.405 0.845 ;
        RECT 945.715 0.515 946.045 0.845 ;
        RECT 944.355 0.515 944.685 0.845 ;
        RECT 942.995 0.515 943.325 0.845 ;
        RECT 941.635 0.515 941.965 0.845 ;
        RECT 940.275 0.515 940.605 0.845 ;
        RECT 938.915 0.515 939.245 0.845 ;
        RECT 937.555 0.515 937.885 0.845 ;
        RECT 936.195 0.515 936.525 0.845 ;
        RECT 934.835 0.515 935.165 0.845 ;
        RECT 933.475 0.515 933.805 0.845 ;
        RECT 932.115 0.515 932.445 0.845 ;
        RECT 930.755 0.515 931.085 0.845 ;
        RECT 929.395 0.515 929.725 0.845 ;
        RECT 928.035 0.515 928.365 0.845 ;
        RECT 926.675 0.515 927.005 0.845 ;
        RECT 925.315 0.515 925.645 0.845 ;
        RECT 923.955 0.515 924.285 0.845 ;
        RECT 922.595 0.515 922.925 0.845 ;
        RECT 921.235 0.515 921.565 0.845 ;
        RECT 919.875 0.515 920.205 0.845 ;
        RECT 918.515 0.515 918.845 0.845 ;
        RECT 917.155 0.515 917.485 0.845 ;
        RECT 915.795 0.515 916.125 0.845 ;
        RECT 914.435 0.515 914.765 0.845 ;
        RECT 913.075 0.515 913.405 0.845 ;
        RECT 911.715 0.515 912.045 0.845 ;
        RECT 910.355 0.515 910.685 0.845 ;
        RECT 908.995 0.515 909.325 0.845 ;
        RECT 907.635 0.515 907.965 0.845 ;
        RECT 906.275 0.515 906.605 0.845 ;
        RECT 904.915 0.515 905.245 0.845 ;
        RECT 903.555 0.515 903.885 0.845 ;
        RECT 902.195 0.515 902.525 0.845 ;
        RECT 900.835 0.515 901.165 0.845 ;
        RECT 899.475 0.515 899.805 0.845 ;
        RECT 898.115 0.515 898.445 0.845 ;
        RECT 896.755 0.515 897.085 0.845 ;
        RECT 895.395 0.515 895.725 0.845 ;
        RECT 894.035 0.515 894.365 0.845 ;
        RECT 892.675 0.515 893.005 0.845 ;
        RECT 891.315 0.515 891.645 0.845 ;
        RECT 889.955 0.515 890.285 0.845 ;
        RECT 888.595 0.515 888.925 0.845 ;
        RECT 887.235 0.515 887.565 0.845 ;
        RECT 885.875 0.515 886.205 0.845 ;
        RECT 884.515 0.515 884.845 0.845 ;
        RECT 883.155 0.515 883.485 0.845 ;
        RECT 881.795 0.515 882.125 0.845 ;
        RECT 880.435 0.515 880.765 0.845 ;
        RECT 879.075 0.515 879.405 0.845 ;
        RECT 877.715 0.515 878.045 0.845 ;
        RECT 876.355 0.515 876.685 0.845 ;
        RECT 874.995 0.515 875.325 0.845 ;
        RECT 873.635 0.515 873.965 0.845 ;
        RECT 872.275 0.515 872.605 0.845 ;
        RECT 870.915 0.515 871.245 0.845 ;
        RECT 869.555 0.515 869.885 0.845 ;
        RECT 868.195 0.515 868.525 0.845 ;
        RECT 866.835 0.515 867.165 0.845 ;
        RECT 865.475 0.515 865.805 0.845 ;
        RECT 864.115 0.515 864.445 0.845 ;
        RECT 862.755 0.515 863.085 0.845 ;
        RECT 861.395 0.515 861.725 0.845 ;
        RECT 860.035 0.515 860.365 0.845 ;
        RECT 858.675 0.515 859.005 0.845 ;
        RECT 857.315 0.515 857.645 0.845 ;
        RECT 855.955 0.515 856.285 0.845 ;
        RECT 854.595 0.515 854.925 0.845 ;
        RECT 853.235 0.515 853.565 0.845 ;
        RECT 851.875 0.515 852.205 0.845 ;
        RECT 850.515 0.515 850.845 0.845 ;
        RECT 849.155 0.515 849.485 0.845 ;
        RECT 847.795 0.515 848.125 0.845 ;
        RECT 846.435 0.515 846.765 0.845 ;
        RECT 845.075 0.515 845.405 0.845 ;
        RECT 843.715 0.515 844.045 0.845 ;
        RECT 842.355 0.515 842.685 0.845 ;
        RECT 840.995 0.515 841.325 0.845 ;
        RECT 839.635 0.515 839.965 0.845 ;
        RECT 838.275 0.515 838.605 0.845 ;
        RECT 836.915 0.515 837.245 0.845 ;
        RECT 835.555 0.515 835.885 0.845 ;
        RECT 834.195 0.515 834.525 0.845 ;
        RECT 832.835 0.515 833.165 0.845 ;
        RECT 831.475 0.515 831.805 0.845 ;
        RECT 830.115 0.515 830.445 0.845 ;
        RECT 828.755 0.515 829.085 0.845 ;
        RECT 827.395 0.515 827.725 0.845 ;
        RECT 826.035 0.515 826.365 0.845 ;
        RECT 824.675 0.515 825.005 0.845 ;
        RECT 823.315 0.515 823.645 0.845 ;
        RECT 821.955 0.515 822.285 0.845 ;
        RECT 820.595 0.515 820.925 0.845 ;
        RECT 819.235 0.515 819.565 0.845 ;
        RECT 817.875 0.515 818.205 0.845 ;
        RECT 816.515 0.515 816.845 0.845 ;
        RECT 815.155 0.515 815.485 0.845 ;
        RECT 813.795 0.515 814.125 0.845 ;
        RECT 812.435 0.515 812.765 0.845 ;
        RECT 811.075 0.515 811.405 0.845 ;
        RECT 809.715 0.515 810.045 0.845 ;
        RECT 808.355 0.515 808.685 0.845 ;
        RECT 806.995 0.515 807.325 0.845 ;
        RECT 805.635 0.515 805.965 0.845 ;
        RECT 804.275 0.515 804.605 0.845 ;
        RECT 802.915 0.515 803.245 0.845 ;
        RECT 801.555 0.515 801.885 0.845 ;
        RECT 800.195 0.515 800.525 0.845 ;
        RECT 798.835 0.515 799.165 0.845 ;
        RECT 797.475 0.515 797.805 0.845 ;
        RECT 796.115 0.515 796.445 0.845 ;
        RECT 794.755 0.515 795.085 0.845 ;
        RECT 793.395 0.515 793.725 0.845 ;
        RECT 792.035 0.515 792.365 0.845 ;
        RECT 790.675 0.515 791.005 0.845 ;
        RECT 789.315 0.515 789.645 0.845 ;
        RECT 787.955 0.515 788.285 0.845 ;
        RECT 786.595 0.515 786.925 0.845 ;
        RECT 785.235 0.515 785.565 0.845 ;
        RECT 783.875 0.515 784.205 0.845 ;
        RECT 782.515 0.515 782.845 0.845 ;
        RECT 781.155 0.515 781.485 0.845 ;
        RECT 779.795 0.515 780.125 0.845 ;
        RECT 778.435 0.515 778.765 0.845 ;
        RECT 777.075 0.515 777.405 0.845 ;
        RECT 775.715 0.515 776.045 0.845 ;
        RECT 774.355 0.515 774.685 0.845 ;
        RECT 772.995 0.515 773.325 0.845 ;
        RECT 771.635 0.515 771.965 0.845 ;
        RECT 770.275 0.515 770.605 0.845 ;
        RECT 768.915 0.515 769.245 0.845 ;
        RECT 767.555 0.515 767.885 0.845 ;
        RECT 766.195 0.515 766.525 0.845 ;
        RECT 764.835 0.515 765.165 0.845 ;
        RECT 763.475 0.515 763.805 0.845 ;
        RECT 762.115 0.515 762.445 0.845 ;
        RECT 760.755 0.515 761.085 0.845 ;
        RECT 759.395 0.515 759.725 0.845 ;
        RECT 758.035 0.515 758.365 0.845 ;
        RECT 756.675 0.515 757.005 0.845 ;
        RECT 755.315 0.515 755.645 0.845 ;
        RECT 753.955 0.515 754.285 0.845 ;
        RECT 752.595 0.515 752.925 0.845 ;
        RECT 751.235 0.515 751.565 0.845 ;
        RECT 749.875 0.515 750.205 0.845 ;
        RECT 748.515 0.515 748.845 0.845 ;
        RECT 747.155 0.515 747.485 0.845 ;
        RECT 745.795 0.515 746.125 0.845 ;
        RECT 744.435 0.515 744.765 0.845 ;
        RECT 743.075 0.515 743.405 0.845 ;
        RECT 741.715 0.515 742.045 0.845 ;
        RECT 740.355 0.515 740.685 0.845 ;
        RECT 738.995 0.515 739.325 0.845 ;
        RECT 737.635 0.515 737.965 0.845 ;
        RECT 736.275 0.515 736.605 0.845 ;
        RECT 734.915 0.515 735.245 0.845 ;
        RECT 733.555 0.515 733.885 0.845 ;
        RECT 732.195 0.515 732.525 0.845 ;
        RECT 730.835 0.515 731.165 0.845 ;
        RECT 729.475 0.515 729.805 0.845 ;
        RECT 728.115 0.515 728.445 0.845 ;
        RECT 726.755 0.515 727.085 0.845 ;
        RECT 725.395 0.515 725.725 0.845 ;
        RECT 724.035 0.515 724.365 0.845 ;
        RECT 722.675 0.515 723.005 0.845 ;
        RECT 721.315 0.515 721.645 0.845 ;
        RECT 719.955 0.515 720.285 0.845 ;
        RECT 718.595 0.515 718.925 0.845 ;
        RECT 717.235 0.515 717.565 0.845 ;
        RECT 715.875 0.515 716.205 0.845 ;
        RECT 714.515 0.515 714.845 0.845 ;
        RECT 713.155 0.515 713.485 0.845 ;
        RECT 711.795 0.515 712.125 0.845 ;
        RECT 710.435 0.515 710.765 0.845 ;
        RECT 709.075 0.515 709.405 0.845 ;
        RECT 707.715 0.515 708.045 0.845 ;
        RECT 706.355 0.515 706.685 0.845 ;
        RECT 704.995 0.515 705.325 0.845 ;
        RECT 703.635 0.515 703.965 0.845 ;
        RECT 702.275 0.515 702.605 0.845 ;
        RECT 700.915 0.515 701.245 0.845 ;
        RECT 699.555 0.515 699.885 0.845 ;
        RECT 698.195 0.515 698.525 0.845 ;
        RECT 696.835 0.515 697.165 0.845 ;
        RECT 695.475 0.515 695.805 0.845 ;
        RECT 694.115 0.515 694.445 0.845 ;
        RECT 692.755 0.515 693.085 0.845 ;
        RECT 691.395 0.515 691.725 0.845 ;
        RECT 690.035 0.515 690.365 0.845 ;
        RECT 688.675 0.515 689.005 0.845 ;
        RECT 687.315 0.515 687.645 0.845 ;
        RECT 685.955 0.515 686.285 0.845 ;
        RECT 684.595 0.515 684.925 0.845 ;
        RECT 683.235 0.515 683.565 0.845 ;
        RECT 681.875 0.515 682.205 0.845 ;
        RECT 680.515 0.515 680.845 0.845 ;
        RECT 679.155 0.515 679.485 0.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -0.845 139.565 -0.515 ;
        RECT 137.875 -0.845 138.205 -0.515 ;
        RECT 136.515 -0.845 136.845 -0.515 ;
        RECT 135.155 -0.845 135.485 -0.515 ;
        RECT 133.795 -0.845 134.125 -0.515 ;
        RECT 132.435 -0.845 132.765 -0.515 ;
        RECT 131.075 -0.845 131.405 -0.515 ;
        RECT 129.715 -0.845 130.045 -0.515 ;
        RECT 128.355 -0.845 128.685 -0.515 ;
        RECT 126.995 -0.845 127.325 -0.515 ;
        RECT 125.635 -0.845 125.965 -0.515 ;
        RECT 124.275 -0.845 124.605 -0.515 ;
        RECT 122.915 -0.845 123.245 -0.515 ;
        RECT 121.555 -0.845 121.885 -0.515 ;
        RECT 120.195 -0.845 120.525 -0.515 ;
        RECT 118.835 -0.845 119.165 -0.515 ;
        RECT 117.475 -0.845 117.805 -0.515 ;
        RECT 116.115 -0.845 116.445 -0.515 ;
        RECT 114.755 -0.845 115.085 -0.515 ;
        RECT 113.395 -0.845 113.725 -0.515 ;
        RECT 112.035 -0.845 112.365 -0.515 ;
        RECT 110.675 -0.845 111.005 -0.515 ;
        RECT 109.315 -0.845 109.645 -0.515 ;
        RECT 107.955 -0.845 108.285 -0.515 ;
        RECT 106.595 -0.845 106.925 -0.515 ;
        RECT 105.235 -0.845 105.565 -0.515 ;
        RECT 103.875 -0.845 104.205 -0.515 ;
        RECT 102.515 -0.845 102.845 -0.515 ;
        RECT 101.155 -0.845 101.485 -0.515 ;
        RECT 99.795 -0.845 100.125 -0.515 ;
        RECT 98.435 -0.845 98.765 -0.515 ;
        RECT 97.075 -0.845 97.405 -0.515 ;
        RECT 95.715 -0.845 96.045 -0.515 ;
        RECT 94.355 -0.845 94.685 -0.515 ;
        RECT 92.995 -0.845 93.325 -0.515 ;
        RECT 91.635 -0.845 91.965 -0.515 ;
        RECT 90.275 -0.845 90.605 -0.515 ;
        RECT 88.915 -0.845 89.245 -0.515 ;
        RECT 87.555 -0.845 87.885 -0.515 ;
        RECT 86.195 -0.845 86.525 -0.515 ;
        RECT 84.835 -0.845 85.165 -0.515 ;
        RECT 83.475 -0.845 83.805 -0.515 ;
        RECT 82.115 -0.845 82.445 -0.515 ;
        RECT 80.755 -0.845 81.085 -0.515 ;
        RECT 79.395 -0.845 79.725 -0.515 ;
        RECT 78.035 -0.845 78.365 -0.515 ;
        RECT 76.675 -0.845 77.005 -0.515 ;
        RECT 75.315 -0.845 75.645 -0.515 ;
        RECT 73.955 -0.845 74.285 -0.515 ;
        RECT 72.595 -0.845 72.925 -0.515 ;
        RECT 71.235 -0.845 71.565 -0.515 ;
        RECT 69.875 -0.845 70.205 -0.515 ;
        RECT 68.515 -0.845 68.845 -0.515 ;
        RECT 67.155 -0.845 67.485 -0.515 ;
        RECT 65.795 -0.845 66.125 -0.515 ;
        RECT 64.435 -0.845 64.765 -0.515 ;
        RECT 63.075 -0.845 63.405 -0.515 ;
        RECT 61.715 -0.845 62.045 -0.515 ;
        RECT 60.355 -0.845 60.685 -0.515 ;
        RECT 58.995 -0.845 59.325 -0.515 ;
        RECT 57.635 -0.845 57.965 -0.515 ;
        RECT 56.275 -0.845 56.605 -0.515 ;
        RECT 54.915 -0.845 55.245 -0.515 ;
        RECT 53.555 -0.845 53.885 -0.515 ;
        RECT 52.195 -0.845 52.525 -0.515 ;
        RECT 50.835 -0.845 51.165 -0.515 ;
        RECT 49.475 -0.845 49.805 -0.515 ;
        RECT 48.115 -0.845 48.445 -0.515 ;
        RECT 46.755 -0.845 47.085 -0.515 ;
        RECT 45.395 -0.845 45.725 -0.515 ;
        RECT 44.035 -0.845 44.365 -0.515 ;
        RECT 42.675 -0.845 43.005 -0.515 ;
        RECT 41.315 -0.845 41.645 -0.515 ;
        RECT 39.955 -0.845 40.285 -0.515 ;
        RECT 38.595 -0.845 38.925 -0.515 ;
        RECT 37.235 -0.845 37.565 -0.515 ;
        RECT 35.875 -0.845 36.205 -0.515 ;
        RECT 34.515 -0.845 34.845 -0.515 ;
        RECT 33.155 -0.845 33.485 -0.515 ;
        RECT 31.795 -0.845 32.125 -0.515 ;
        RECT 30.435 -0.845 30.765 -0.515 ;
        RECT 29.075 -0.845 29.405 -0.515 ;
        RECT 27.715 -0.845 28.045 -0.515 ;
        RECT 26.355 -0.845 26.685 -0.515 ;
        RECT 24.995 -0.845 25.325 -0.515 ;
        RECT 23.635 -0.845 23.965 -0.515 ;
        RECT 22.275 -0.845 22.605 -0.515 ;
        RECT 20.915 -0.845 21.245 -0.515 ;
        RECT 19.555 -0.845 19.885 -0.515 ;
        RECT 18.195 -0.845 18.525 -0.515 ;
        RECT 16.835 -0.845 17.165 -0.515 ;
        RECT 15.475 -0.845 15.805 -0.515 ;
        RECT 14.115 -0.845 14.445 -0.515 ;
        RECT 12.755 -0.845 13.085 -0.515 ;
        RECT 11.395 -0.845 11.725 -0.515 ;
        RECT 10.035 -0.845 10.365 -0.515 ;
        RECT 8.675 -0.845 9.005 -0.515 ;
        RECT 7.315 -0.845 7.645 -0.515 ;
        RECT 5.955 -0.845 6.285 -0.515 ;
        RECT 4.595 -0.845 4.925 -0.515 ;
        RECT 3.235 -0.845 3.565 -0.515 ;
        RECT 1.875 -0.845 2.205 -0.515 ;
        RECT 0.515 -0.845 0.845 -0.515 ;
        RECT -0.845 -0.845 -0.515 -0.515 ;
        RECT 677.795 -0.845 678.125 -0.515 ;
        RECT -1.52 -0.84 678.125 -0.52 ;
        RECT 676.435 -0.845 676.765 -0.515 ;
        RECT 675.075 -0.845 675.405 -0.515 ;
        RECT 673.715 -0.845 674.045 -0.515 ;
        RECT 672.355 -0.845 672.685 -0.515 ;
        RECT 670.995 -0.845 671.325 -0.515 ;
        RECT 669.635 -0.845 669.965 -0.515 ;
        RECT 668.275 -0.845 668.605 -0.515 ;
        RECT 666.915 -0.845 667.245 -0.515 ;
        RECT 665.555 -0.845 665.885 -0.515 ;
        RECT 664.195 -0.845 664.525 -0.515 ;
        RECT 662.835 -0.845 663.165 -0.515 ;
        RECT 661.475 -0.845 661.805 -0.515 ;
        RECT 660.115 -0.845 660.445 -0.515 ;
        RECT 658.755 -0.845 659.085 -0.515 ;
        RECT 657.395 -0.845 657.725 -0.515 ;
        RECT 656.035 -0.845 656.365 -0.515 ;
        RECT 654.675 -0.845 655.005 -0.515 ;
        RECT 653.315 -0.845 653.645 -0.515 ;
        RECT 651.955 -0.845 652.285 -0.515 ;
        RECT 650.595 -0.845 650.925 -0.515 ;
        RECT 649.235 -0.845 649.565 -0.515 ;
        RECT 647.875 -0.845 648.205 -0.515 ;
        RECT 646.515 -0.845 646.845 -0.515 ;
        RECT 645.155 -0.845 645.485 -0.515 ;
        RECT 643.795 -0.845 644.125 -0.515 ;
        RECT 642.435 -0.845 642.765 -0.515 ;
        RECT 641.075 -0.845 641.405 -0.515 ;
        RECT 639.715 -0.845 640.045 -0.515 ;
        RECT 638.355 -0.845 638.685 -0.515 ;
        RECT 636.995 -0.845 637.325 -0.515 ;
        RECT 635.635 -0.845 635.965 -0.515 ;
        RECT 634.275 -0.845 634.605 -0.515 ;
        RECT 632.915 -0.845 633.245 -0.515 ;
        RECT 631.555 -0.845 631.885 -0.515 ;
        RECT 630.195 -0.845 630.525 -0.515 ;
        RECT 628.835 -0.845 629.165 -0.515 ;
        RECT 627.475 -0.845 627.805 -0.515 ;
        RECT 626.115 -0.845 626.445 -0.515 ;
        RECT 624.755 -0.845 625.085 -0.515 ;
        RECT 623.395 -0.845 623.725 -0.515 ;
        RECT 622.035 -0.845 622.365 -0.515 ;
        RECT 620.675 -0.845 621.005 -0.515 ;
        RECT 619.315 -0.845 619.645 -0.515 ;
        RECT 617.955 -0.845 618.285 -0.515 ;
        RECT 616.595 -0.845 616.925 -0.515 ;
        RECT 615.235 -0.845 615.565 -0.515 ;
        RECT 613.875 -0.845 614.205 -0.515 ;
        RECT 612.515 -0.845 612.845 -0.515 ;
        RECT 611.155 -0.845 611.485 -0.515 ;
        RECT 609.795 -0.845 610.125 -0.515 ;
        RECT 608.435 -0.845 608.765 -0.515 ;
        RECT 607.075 -0.845 607.405 -0.515 ;
        RECT 605.715 -0.845 606.045 -0.515 ;
        RECT 604.355 -0.845 604.685 -0.515 ;
        RECT 602.995 -0.845 603.325 -0.515 ;
        RECT 601.635 -0.845 601.965 -0.515 ;
        RECT 600.275 -0.845 600.605 -0.515 ;
        RECT 598.915 -0.845 599.245 -0.515 ;
        RECT 597.555 -0.845 597.885 -0.515 ;
        RECT 596.195 -0.845 596.525 -0.515 ;
        RECT 594.835 -0.845 595.165 -0.515 ;
        RECT 593.475 -0.845 593.805 -0.515 ;
        RECT 592.115 -0.845 592.445 -0.515 ;
        RECT 590.755 -0.845 591.085 -0.515 ;
        RECT 589.395 -0.845 589.725 -0.515 ;
        RECT 588.035 -0.845 588.365 -0.515 ;
        RECT 586.675 -0.845 587.005 -0.515 ;
        RECT 585.315 -0.845 585.645 -0.515 ;
        RECT 583.955 -0.845 584.285 -0.515 ;
        RECT 582.595 -0.845 582.925 -0.515 ;
        RECT 581.235 -0.845 581.565 -0.515 ;
        RECT 579.875 -0.845 580.205 -0.515 ;
        RECT 578.515 -0.845 578.845 -0.515 ;
        RECT 577.155 -0.845 577.485 -0.515 ;
        RECT 575.795 -0.845 576.125 -0.515 ;
        RECT 574.435 -0.845 574.765 -0.515 ;
        RECT 573.075 -0.845 573.405 -0.515 ;
        RECT 571.715 -0.845 572.045 -0.515 ;
        RECT 570.355 -0.845 570.685 -0.515 ;
        RECT 568.995 -0.845 569.325 -0.515 ;
        RECT 567.635 -0.845 567.965 -0.515 ;
        RECT 566.275 -0.845 566.605 -0.515 ;
        RECT 564.915 -0.845 565.245 -0.515 ;
        RECT 563.555 -0.845 563.885 -0.515 ;
        RECT 562.195 -0.845 562.525 -0.515 ;
        RECT 560.835 -0.845 561.165 -0.515 ;
        RECT 559.475 -0.845 559.805 -0.515 ;
        RECT 558.115 -0.845 558.445 -0.515 ;
        RECT 556.755 -0.845 557.085 -0.515 ;
        RECT 555.395 -0.845 555.725 -0.515 ;
        RECT 554.035 -0.845 554.365 -0.515 ;
        RECT 552.675 -0.845 553.005 -0.515 ;
        RECT 551.315 -0.845 551.645 -0.515 ;
        RECT 549.955 -0.845 550.285 -0.515 ;
        RECT 548.595 -0.845 548.925 -0.515 ;
        RECT 547.235 -0.845 547.565 -0.515 ;
        RECT 545.875 -0.845 546.205 -0.515 ;
        RECT 544.515 -0.845 544.845 -0.515 ;
        RECT 543.155 -0.845 543.485 -0.515 ;
        RECT 541.795 -0.845 542.125 -0.515 ;
        RECT 540.435 -0.845 540.765 -0.515 ;
        RECT 539.075 -0.845 539.405 -0.515 ;
        RECT 537.715 -0.845 538.045 -0.515 ;
        RECT 536.355 -0.845 536.685 -0.515 ;
        RECT 534.995 -0.845 535.325 -0.515 ;
        RECT 533.635 -0.845 533.965 -0.515 ;
        RECT 532.275 -0.845 532.605 -0.515 ;
        RECT 530.915 -0.845 531.245 -0.515 ;
        RECT 529.555 -0.845 529.885 -0.515 ;
        RECT 528.195 -0.845 528.525 -0.515 ;
        RECT 526.835 -0.845 527.165 -0.515 ;
        RECT 525.475 -0.845 525.805 -0.515 ;
        RECT 524.115 -0.845 524.445 -0.515 ;
        RECT 522.755 -0.845 523.085 -0.515 ;
        RECT 521.395 -0.845 521.725 -0.515 ;
        RECT 520.035 -0.845 520.365 -0.515 ;
        RECT 518.675 -0.845 519.005 -0.515 ;
        RECT 517.315 -0.845 517.645 -0.515 ;
        RECT 515.955 -0.845 516.285 -0.515 ;
        RECT 514.595 -0.845 514.925 -0.515 ;
        RECT 513.235 -0.845 513.565 -0.515 ;
        RECT 511.875 -0.845 512.205 -0.515 ;
        RECT 510.515 -0.845 510.845 -0.515 ;
        RECT 509.155 -0.845 509.485 -0.515 ;
        RECT 507.795 -0.845 508.125 -0.515 ;
        RECT 506.435 -0.845 506.765 -0.515 ;
        RECT 505.075 -0.845 505.405 -0.515 ;
        RECT 503.715 -0.845 504.045 -0.515 ;
        RECT 502.355 -0.845 502.685 -0.515 ;
        RECT 500.995 -0.845 501.325 -0.515 ;
        RECT 499.635 -0.845 499.965 -0.515 ;
        RECT 498.275 -0.845 498.605 -0.515 ;
        RECT 496.915 -0.845 497.245 -0.515 ;
        RECT 495.555 -0.845 495.885 -0.515 ;
        RECT 494.195 -0.845 494.525 -0.515 ;
        RECT 492.835 -0.845 493.165 -0.515 ;
        RECT 491.475 -0.845 491.805 -0.515 ;
        RECT 490.115 -0.845 490.445 -0.515 ;
        RECT 488.755 -0.845 489.085 -0.515 ;
        RECT 487.395 -0.845 487.725 -0.515 ;
        RECT 486.035 -0.845 486.365 -0.515 ;
        RECT 484.675 -0.845 485.005 -0.515 ;
        RECT 483.315 -0.845 483.645 -0.515 ;
        RECT 481.955 -0.845 482.285 -0.515 ;
        RECT 480.595 -0.845 480.925 -0.515 ;
        RECT 479.235 -0.845 479.565 -0.515 ;
        RECT 477.875 -0.845 478.205 -0.515 ;
        RECT 476.515 -0.845 476.845 -0.515 ;
        RECT 475.155 -0.845 475.485 -0.515 ;
        RECT 473.795 -0.845 474.125 -0.515 ;
        RECT 472.435 -0.845 472.765 -0.515 ;
        RECT 471.075 -0.845 471.405 -0.515 ;
        RECT 469.715 -0.845 470.045 -0.515 ;
        RECT 468.355 -0.845 468.685 -0.515 ;
        RECT 466.995 -0.845 467.325 -0.515 ;
        RECT 465.635 -0.845 465.965 -0.515 ;
        RECT 464.275 -0.845 464.605 -0.515 ;
        RECT 462.915 -0.845 463.245 -0.515 ;
        RECT 461.555 -0.845 461.885 -0.515 ;
        RECT 460.195 -0.845 460.525 -0.515 ;
        RECT 458.835 -0.845 459.165 -0.515 ;
        RECT 457.475 -0.845 457.805 -0.515 ;
        RECT 456.115 -0.845 456.445 -0.515 ;
        RECT 454.755 -0.845 455.085 -0.515 ;
        RECT 453.395 -0.845 453.725 -0.515 ;
        RECT 452.035 -0.845 452.365 -0.515 ;
        RECT 450.675 -0.845 451.005 -0.515 ;
        RECT 449.315 -0.845 449.645 -0.515 ;
        RECT 447.955 -0.845 448.285 -0.515 ;
        RECT 446.595 -0.845 446.925 -0.515 ;
        RECT 445.235 -0.845 445.565 -0.515 ;
        RECT 443.875 -0.845 444.205 -0.515 ;
        RECT 442.515 -0.845 442.845 -0.515 ;
        RECT 441.155 -0.845 441.485 -0.515 ;
        RECT 439.795 -0.845 440.125 -0.515 ;
        RECT 438.435 -0.845 438.765 -0.515 ;
        RECT 437.075 -0.845 437.405 -0.515 ;
        RECT 435.715 -0.845 436.045 -0.515 ;
        RECT 434.355 -0.845 434.685 -0.515 ;
        RECT 432.995 -0.845 433.325 -0.515 ;
        RECT 431.635 -0.845 431.965 -0.515 ;
        RECT 430.275 -0.845 430.605 -0.515 ;
        RECT 428.915 -0.845 429.245 -0.515 ;
        RECT 427.555 -0.845 427.885 -0.515 ;
        RECT 426.195 -0.845 426.525 -0.515 ;
        RECT 424.835 -0.845 425.165 -0.515 ;
        RECT 423.475 -0.845 423.805 -0.515 ;
        RECT 422.115 -0.845 422.445 -0.515 ;
        RECT 420.755 -0.845 421.085 -0.515 ;
        RECT 419.395 -0.845 419.725 -0.515 ;
        RECT 418.035 -0.845 418.365 -0.515 ;
        RECT 416.675 -0.845 417.005 -0.515 ;
        RECT 415.315 -0.845 415.645 -0.515 ;
        RECT 413.955 -0.845 414.285 -0.515 ;
        RECT 412.595 -0.845 412.925 -0.515 ;
        RECT 411.235 -0.845 411.565 -0.515 ;
        RECT 409.875 -0.845 410.205 -0.515 ;
        RECT 408.515 -0.845 408.845 -0.515 ;
        RECT 407.155 -0.845 407.485 -0.515 ;
        RECT 405.795 -0.845 406.125 -0.515 ;
        RECT 404.435 -0.845 404.765 -0.515 ;
        RECT 403.075 -0.845 403.405 -0.515 ;
        RECT 401.715 -0.845 402.045 -0.515 ;
        RECT 400.355 -0.845 400.685 -0.515 ;
        RECT 398.995 -0.845 399.325 -0.515 ;
        RECT 397.635 -0.845 397.965 -0.515 ;
        RECT 396.275 -0.845 396.605 -0.515 ;
        RECT 394.915 -0.845 395.245 -0.515 ;
        RECT 393.555 -0.845 393.885 -0.515 ;
        RECT 392.195 -0.845 392.525 -0.515 ;
        RECT 390.835 -0.845 391.165 -0.515 ;
        RECT 389.475 -0.845 389.805 -0.515 ;
        RECT 388.115 -0.845 388.445 -0.515 ;
        RECT 386.755 -0.845 387.085 -0.515 ;
        RECT 385.395 -0.845 385.725 -0.515 ;
        RECT 384.035 -0.845 384.365 -0.515 ;
        RECT 382.675 -0.845 383.005 -0.515 ;
        RECT 381.315 -0.845 381.645 -0.515 ;
        RECT 379.955 -0.845 380.285 -0.515 ;
        RECT 378.595 -0.845 378.925 -0.515 ;
        RECT 377.235 -0.845 377.565 -0.515 ;
        RECT 375.875 -0.845 376.205 -0.515 ;
        RECT 374.515 -0.845 374.845 -0.515 ;
        RECT 373.155 -0.845 373.485 -0.515 ;
        RECT 371.795 -0.845 372.125 -0.515 ;
        RECT 370.435 -0.845 370.765 -0.515 ;
        RECT 369.075 -0.845 369.405 -0.515 ;
        RECT 367.715 -0.845 368.045 -0.515 ;
        RECT 366.355 -0.845 366.685 -0.515 ;
        RECT 364.995 -0.845 365.325 -0.515 ;
        RECT 363.635 -0.845 363.965 -0.515 ;
        RECT 362.275 -0.845 362.605 -0.515 ;
        RECT 360.915 -0.845 361.245 -0.515 ;
        RECT 359.555 -0.845 359.885 -0.515 ;
        RECT 358.195 -0.845 358.525 -0.515 ;
        RECT 356.835 -0.845 357.165 -0.515 ;
        RECT 355.475 -0.845 355.805 -0.515 ;
        RECT 354.115 -0.845 354.445 -0.515 ;
        RECT 352.755 -0.845 353.085 -0.515 ;
        RECT 351.395 -0.845 351.725 -0.515 ;
        RECT 350.035 -0.845 350.365 -0.515 ;
        RECT 348.675 -0.845 349.005 -0.515 ;
        RECT 347.315 -0.845 347.645 -0.515 ;
        RECT 345.955 -0.845 346.285 -0.515 ;
        RECT 344.595 -0.845 344.925 -0.515 ;
        RECT 343.235 -0.845 343.565 -0.515 ;
        RECT 341.875 -0.845 342.205 -0.515 ;
        RECT 340.515 -0.845 340.845 -0.515 ;
        RECT 339.155 -0.845 339.485 -0.515 ;
        RECT 337.795 -0.845 338.125 -0.515 ;
        RECT 336.435 -0.845 336.765 -0.515 ;
        RECT 335.075 -0.845 335.405 -0.515 ;
        RECT 333.715 -0.845 334.045 -0.515 ;
        RECT 332.355 -0.845 332.685 -0.515 ;
        RECT 330.995 -0.845 331.325 -0.515 ;
        RECT 329.635 -0.845 329.965 -0.515 ;
        RECT 328.275 -0.845 328.605 -0.515 ;
        RECT 326.915 -0.845 327.245 -0.515 ;
        RECT 325.555 -0.845 325.885 -0.515 ;
        RECT 324.195 -0.845 324.525 -0.515 ;
        RECT 322.835 -0.845 323.165 -0.515 ;
        RECT 321.475 -0.845 321.805 -0.515 ;
        RECT 320.115 -0.845 320.445 -0.515 ;
        RECT 318.755 -0.845 319.085 -0.515 ;
        RECT 317.395 -0.845 317.725 -0.515 ;
        RECT 316.035 -0.845 316.365 -0.515 ;
        RECT 314.675 -0.845 315.005 -0.515 ;
        RECT 313.315 -0.845 313.645 -0.515 ;
        RECT 311.955 -0.845 312.285 -0.515 ;
        RECT 310.595 -0.845 310.925 -0.515 ;
        RECT 309.235 -0.845 309.565 -0.515 ;
        RECT 307.875 -0.845 308.205 -0.515 ;
        RECT 306.515 -0.845 306.845 -0.515 ;
        RECT 305.155 -0.845 305.485 -0.515 ;
        RECT 303.795 -0.845 304.125 -0.515 ;
        RECT 302.435 -0.845 302.765 -0.515 ;
        RECT 301.075 -0.845 301.405 -0.515 ;
        RECT 299.715 -0.845 300.045 -0.515 ;
        RECT 298.355 -0.845 298.685 -0.515 ;
        RECT 296.995 -0.845 297.325 -0.515 ;
        RECT 295.635 -0.845 295.965 -0.515 ;
        RECT 294.275 -0.845 294.605 -0.515 ;
        RECT 292.915 -0.845 293.245 -0.515 ;
        RECT 291.555 -0.845 291.885 -0.515 ;
        RECT 290.195 -0.845 290.525 -0.515 ;
        RECT 288.835 -0.845 289.165 -0.515 ;
        RECT 287.475 -0.845 287.805 -0.515 ;
        RECT 286.115 -0.845 286.445 -0.515 ;
        RECT 284.755 -0.845 285.085 -0.515 ;
        RECT 283.395 -0.845 283.725 -0.515 ;
        RECT 282.035 -0.845 282.365 -0.515 ;
        RECT 280.675 -0.845 281.005 -0.515 ;
        RECT 279.315 -0.845 279.645 -0.515 ;
        RECT 277.955 -0.845 278.285 -0.515 ;
        RECT 276.595 -0.845 276.925 -0.515 ;
        RECT 275.235 -0.845 275.565 -0.515 ;
        RECT 273.875 -0.845 274.205 -0.515 ;
        RECT 272.515 -0.845 272.845 -0.515 ;
        RECT 271.155 -0.845 271.485 -0.515 ;
        RECT 269.795 -0.845 270.125 -0.515 ;
        RECT 268.435 -0.845 268.765 -0.515 ;
        RECT 267.075 -0.845 267.405 -0.515 ;
        RECT 265.715 -0.845 266.045 -0.515 ;
        RECT 264.355 -0.845 264.685 -0.515 ;
        RECT 262.995 -0.845 263.325 -0.515 ;
        RECT 261.635 -0.845 261.965 -0.515 ;
        RECT 260.275 -0.845 260.605 -0.515 ;
        RECT 258.915 -0.845 259.245 -0.515 ;
        RECT 257.555 -0.845 257.885 -0.515 ;
        RECT 256.195 -0.845 256.525 -0.515 ;
        RECT 254.835 -0.845 255.165 -0.515 ;
        RECT 253.475 -0.845 253.805 -0.515 ;
        RECT 252.115 -0.845 252.445 -0.515 ;
        RECT 250.755 -0.845 251.085 -0.515 ;
        RECT 249.395 -0.845 249.725 -0.515 ;
        RECT 248.035 -0.845 248.365 -0.515 ;
        RECT 246.675 -0.845 247.005 -0.515 ;
        RECT 245.315 -0.845 245.645 -0.515 ;
        RECT 243.955 -0.845 244.285 -0.515 ;
        RECT 242.595 -0.845 242.925 -0.515 ;
        RECT 241.235 -0.845 241.565 -0.515 ;
        RECT 239.875 -0.845 240.205 -0.515 ;
        RECT 238.515 -0.845 238.845 -0.515 ;
        RECT 237.155 -0.845 237.485 -0.515 ;
        RECT 235.795 -0.845 236.125 -0.515 ;
        RECT 234.435 -0.845 234.765 -0.515 ;
        RECT 233.075 -0.845 233.405 -0.515 ;
        RECT 231.715 -0.845 232.045 -0.515 ;
        RECT 230.355 -0.845 230.685 -0.515 ;
        RECT 228.995 -0.845 229.325 -0.515 ;
        RECT 227.635 -0.845 227.965 -0.515 ;
        RECT 226.275 -0.845 226.605 -0.515 ;
        RECT 224.915 -0.845 225.245 -0.515 ;
        RECT 223.555 -0.845 223.885 -0.515 ;
        RECT 222.195 -0.845 222.525 -0.515 ;
        RECT 220.835 -0.845 221.165 -0.515 ;
        RECT 219.475 -0.845 219.805 -0.515 ;
        RECT 218.115 -0.845 218.445 -0.515 ;
        RECT 216.755 -0.845 217.085 -0.515 ;
        RECT 215.395 -0.845 215.725 -0.515 ;
        RECT 214.035 -0.845 214.365 -0.515 ;
        RECT 212.675 -0.845 213.005 -0.515 ;
        RECT 211.315 -0.845 211.645 -0.515 ;
        RECT 209.955 -0.845 210.285 -0.515 ;
        RECT 208.595 -0.845 208.925 -0.515 ;
        RECT 207.235 -0.845 207.565 -0.515 ;
        RECT 205.875 -0.845 206.205 -0.515 ;
        RECT 204.515 -0.845 204.845 -0.515 ;
        RECT 203.155 -0.845 203.485 -0.515 ;
        RECT 201.795 -0.845 202.125 -0.515 ;
        RECT 200.435 -0.845 200.765 -0.515 ;
        RECT 199.075 -0.845 199.405 -0.515 ;
        RECT 197.715 -0.845 198.045 -0.515 ;
        RECT 196.355 -0.845 196.685 -0.515 ;
        RECT 194.995 -0.845 195.325 -0.515 ;
        RECT 193.635 -0.845 193.965 -0.515 ;
        RECT 192.275 -0.845 192.605 -0.515 ;
        RECT 190.915 -0.845 191.245 -0.515 ;
        RECT 189.555 -0.845 189.885 -0.515 ;
        RECT 188.195 -0.845 188.525 -0.515 ;
        RECT 186.835 -0.845 187.165 -0.515 ;
        RECT 185.475 -0.845 185.805 -0.515 ;
        RECT 184.115 -0.845 184.445 -0.515 ;
        RECT 182.755 -0.845 183.085 -0.515 ;
        RECT 181.395 -0.845 181.725 -0.515 ;
        RECT 180.035 -0.845 180.365 -0.515 ;
        RECT 178.675 -0.845 179.005 -0.515 ;
        RECT 177.315 -0.845 177.645 -0.515 ;
        RECT 175.955 -0.845 176.285 -0.515 ;
        RECT 174.595 -0.845 174.925 -0.515 ;
        RECT 173.235 -0.845 173.565 -0.515 ;
        RECT 171.875 -0.845 172.205 -0.515 ;
        RECT 170.515 -0.845 170.845 -0.515 ;
        RECT 169.155 -0.845 169.485 -0.515 ;
        RECT 167.795 -0.845 168.125 -0.515 ;
        RECT 166.435 -0.845 166.765 -0.515 ;
        RECT 165.075 -0.845 165.405 -0.515 ;
        RECT 163.715 -0.845 164.045 -0.515 ;
        RECT 162.355 -0.845 162.685 -0.515 ;
        RECT 160.995 -0.845 161.325 -0.515 ;
        RECT 159.635 -0.845 159.965 -0.515 ;
        RECT 158.275 -0.845 158.605 -0.515 ;
        RECT 156.915 -0.845 157.245 -0.515 ;
        RECT 155.555 -0.845 155.885 -0.515 ;
        RECT 154.195 -0.845 154.525 -0.515 ;
        RECT 152.835 -0.845 153.165 -0.515 ;
        RECT 151.475 -0.845 151.805 -0.515 ;
        RECT 150.115 -0.845 150.445 -0.515 ;
        RECT 148.755 -0.845 149.085 -0.515 ;
        RECT 147.395 -0.845 147.725 -0.515 ;
        RECT 146.035 -0.845 146.365 -0.515 ;
        RECT 144.675 -0.845 145.005 -0.515 ;
        RECT 143.315 -0.845 143.645 -0.515 ;
        RECT 141.955 -0.845 142.285 -0.515 ;
        RECT 140.595 -0.845 140.925 -0.515 ;
        RECT 678.125 -0.84 954.88 -0.52 ;
        RECT 953.875 -0.845 954.205 -0.515 ;
        RECT 952.515 -0.845 952.845 -0.515 ;
        RECT 951.155 -0.845 951.485 -0.515 ;
        RECT 949.795 -0.845 950.125 -0.515 ;
        RECT 948.435 -0.845 948.765 -0.515 ;
        RECT 947.075 -0.845 947.405 -0.515 ;
        RECT 945.715 -0.845 946.045 -0.515 ;
        RECT 944.355 -0.845 944.685 -0.515 ;
        RECT 942.995 -0.845 943.325 -0.515 ;
        RECT 941.635 -0.845 941.965 -0.515 ;
        RECT 940.275 -0.845 940.605 -0.515 ;
        RECT 938.915 -0.845 939.245 -0.515 ;
        RECT 937.555 -0.845 937.885 -0.515 ;
        RECT 936.195 -0.845 936.525 -0.515 ;
        RECT 934.835 -0.845 935.165 -0.515 ;
        RECT 933.475 -0.845 933.805 -0.515 ;
        RECT 932.115 -0.845 932.445 -0.515 ;
        RECT 930.755 -0.845 931.085 -0.515 ;
        RECT 929.395 -0.845 929.725 -0.515 ;
        RECT 928.035 -0.845 928.365 -0.515 ;
        RECT 926.675 -0.845 927.005 -0.515 ;
        RECT 925.315 -0.845 925.645 -0.515 ;
        RECT 923.955 -0.845 924.285 -0.515 ;
        RECT 922.595 -0.845 922.925 -0.515 ;
        RECT 921.235 -0.845 921.565 -0.515 ;
        RECT 919.875 -0.845 920.205 -0.515 ;
        RECT 918.515 -0.845 918.845 -0.515 ;
        RECT 917.155 -0.845 917.485 -0.515 ;
        RECT 915.795 -0.845 916.125 -0.515 ;
        RECT 914.435 -0.845 914.765 -0.515 ;
        RECT 913.075 -0.845 913.405 -0.515 ;
        RECT 911.715 -0.845 912.045 -0.515 ;
        RECT 910.355 -0.845 910.685 -0.515 ;
        RECT 908.995 -0.845 909.325 -0.515 ;
        RECT 907.635 -0.845 907.965 -0.515 ;
        RECT 906.275 -0.845 906.605 -0.515 ;
        RECT 904.915 -0.845 905.245 -0.515 ;
        RECT 903.555 -0.845 903.885 -0.515 ;
        RECT 902.195 -0.845 902.525 -0.515 ;
        RECT 900.835 -0.845 901.165 -0.515 ;
        RECT 899.475 -0.845 899.805 -0.515 ;
        RECT 898.115 -0.845 898.445 -0.515 ;
        RECT 896.755 -0.845 897.085 -0.515 ;
        RECT 895.395 -0.845 895.725 -0.515 ;
        RECT 894.035 -0.845 894.365 -0.515 ;
        RECT 892.675 -0.845 893.005 -0.515 ;
        RECT 891.315 -0.845 891.645 -0.515 ;
        RECT 889.955 -0.845 890.285 -0.515 ;
        RECT 888.595 -0.845 888.925 -0.515 ;
        RECT 887.235 -0.845 887.565 -0.515 ;
        RECT 885.875 -0.845 886.205 -0.515 ;
        RECT 884.515 -0.845 884.845 -0.515 ;
        RECT 883.155 -0.845 883.485 -0.515 ;
        RECT 881.795 -0.845 882.125 -0.515 ;
        RECT 880.435 -0.845 880.765 -0.515 ;
        RECT 879.075 -0.845 879.405 -0.515 ;
        RECT 877.715 -0.845 878.045 -0.515 ;
        RECT 876.355 -0.845 876.685 -0.515 ;
        RECT 874.995 -0.845 875.325 -0.515 ;
        RECT 873.635 -0.845 873.965 -0.515 ;
        RECT 872.275 -0.845 872.605 -0.515 ;
        RECT 870.915 -0.845 871.245 -0.515 ;
        RECT 869.555 -0.845 869.885 -0.515 ;
        RECT 868.195 -0.845 868.525 -0.515 ;
        RECT 866.835 -0.845 867.165 -0.515 ;
        RECT 865.475 -0.845 865.805 -0.515 ;
        RECT 864.115 -0.845 864.445 -0.515 ;
        RECT 862.755 -0.845 863.085 -0.515 ;
        RECT 861.395 -0.845 861.725 -0.515 ;
        RECT 860.035 -0.845 860.365 -0.515 ;
        RECT 858.675 -0.845 859.005 -0.515 ;
        RECT 857.315 -0.845 857.645 -0.515 ;
        RECT 855.955 -0.845 856.285 -0.515 ;
        RECT 854.595 -0.845 854.925 -0.515 ;
        RECT 853.235 -0.845 853.565 -0.515 ;
        RECT 851.875 -0.845 852.205 -0.515 ;
        RECT 850.515 -0.845 850.845 -0.515 ;
        RECT 849.155 -0.845 849.485 -0.515 ;
        RECT 847.795 -0.845 848.125 -0.515 ;
        RECT 846.435 -0.845 846.765 -0.515 ;
        RECT 845.075 -0.845 845.405 -0.515 ;
        RECT 843.715 -0.845 844.045 -0.515 ;
        RECT 842.355 -0.845 842.685 -0.515 ;
        RECT 840.995 -0.845 841.325 -0.515 ;
        RECT 839.635 -0.845 839.965 -0.515 ;
        RECT 838.275 -0.845 838.605 -0.515 ;
        RECT 836.915 -0.845 837.245 -0.515 ;
        RECT 835.555 -0.845 835.885 -0.515 ;
        RECT 834.195 -0.845 834.525 -0.515 ;
        RECT 832.835 -0.845 833.165 -0.515 ;
        RECT 831.475 -0.845 831.805 -0.515 ;
        RECT 830.115 -0.845 830.445 -0.515 ;
        RECT 828.755 -0.845 829.085 -0.515 ;
        RECT 827.395 -0.845 827.725 -0.515 ;
        RECT 826.035 -0.845 826.365 -0.515 ;
        RECT 824.675 -0.845 825.005 -0.515 ;
        RECT 823.315 -0.845 823.645 -0.515 ;
        RECT 821.955 -0.845 822.285 -0.515 ;
        RECT 820.595 -0.845 820.925 -0.515 ;
        RECT 819.235 -0.845 819.565 -0.515 ;
        RECT 817.875 -0.845 818.205 -0.515 ;
        RECT 816.515 -0.845 816.845 -0.515 ;
        RECT 815.155 -0.845 815.485 -0.515 ;
        RECT 813.795 -0.845 814.125 -0.515 ;
        RECT 812.435 -0.845 812.765 -0.515 ;
        RECT 811.075 -0.845 811.405 -0.515 ;
        RECT 809.715 -0.845 810.045 -0.515 ;
        RECT 808.355 -0.845 808.685 -0.515 ;
        RECT 806.995 -0.845 807.325 -0.515 ;
        RECT 805.635 -0.845 805.965 -0.515 ;
        RECT 804.275 -0.845 804.605 -0.515 ;
        RECT 802.915 -0.845 803.245 -0.515 ;
        RECT 801.555 -0.845 801.885 -0.515 ;
        RECT 800.195 -0.845 800.525 -0.515 ;
        RECT 798.835 -0.845 799.165 -0.515 ;
        RECT 797.475 -0.845 797.805 -0.515 ;
        RECT 796.115 -0.845 796.445 -0.515 ;
        RECT 794.755 -0.845 795.085 -0.515 ;
        RECT 793.395 -0.845 793.725 -0.515 ;
        RECT 792.035 -0.845 792.365 -0.515 ;
        RECT 790.675 -0.845 791.005 -0.515 ;
        RECT 789.315 -0.845 789.645 -0.515 ;
        RECT 787.955 -0.845 788.285 -0.515 ;
        RECT 786.595 -0.845 786.925 -0.515 ;
        RECT 785.235 -0.845 785.565 -0.515 ;
        RECT 783.875 -0.845 784.205 -0.515 ;
        RECT 782.515 -0.845 782.845 -0.515 ;
        RECT 781.155 -0.845 781.485 -0.515 ;
        RECT 779.795 -0.845 780.125 -0.515 ;
        RECT 778.435 -0.845 778.765 -0.515 ;
        RECT 777.075 -0.845 777.405 -0.515 ;
        RECT 775.715 -0.845 776.045 -0.515 ;
        RECT 774.355 -0.845 774.685 -0.515 ;
        RECT 772.995 -0.845 773.325 -0.515 ;
        RECT 771.635 -0.845 771.965 -0.515 ;
        RECT 770.275 -0.845 770.605 -0.515 ;
        RECT 768.915 -0.845 769.245 -0.515 ;
        RECT 767.555 -0.845 767.885 -0.515 ;
        RECT 766.195 -0.845 766.525 -0.515 ;
        RECT 764.835 -0.845 765.165 -0.515 ;
        RECT 763.475 -0.845 763.805 -0.515 ;
        RECT 762.115 -0.845 762.445 -0.515 ;
        RECT 760.755 -0.845 761.085 -0.515 ;
        RECT 759.395 -0.845 759.725 -0.515 ;
        RECT 758.035 -0.845 758.365 -0.515 ;
        RECT 756.675 -0.845 757.005 -0.515 ;
        RECT 755.315 -0.845 755.645 -0.515 ;
        RECT 753.955 -0.845 754.285 -0.515 ;
        RECT 752.595 -0.845 752.925 -0.515 ;
        RECT 751.235 -0.845 751.565 -0.515 ;
        RECT 749.875 -0.845 750.205 -0.515 ;
        RECT 748.515 -0.845 748.845 -0.515 ;
        RECT 747.155 -0.845 747.485 -0.515 ;
        RECT 745.795 -0.845 746.125 -0.515 ;
        RECT 744.435 -0.845 744.765 -0.515 ;
        RECT 743.075 -0.845 743.405 -0.515 ;
        RECT 741.715 -0.845 742.045 -0.515 ;
        RECT 740.355 -0.845 740.685 -0.515 ;
        RECT 738.995 -0.845 739.325 -0.515 ;
        RECT 737.635 -0.845 737.965 -0.515 ;
        RECT 736.275 -0.845 736.605 -0.515 ;
        RECT 734.915 -0.845 735.245 -0.515 ;
        RECT 733.555 -0.845 733.885 -0.515 ;
        RECT 732.195 -0.845 732.525 -0.515 ;
        RECT 730.835 -0.845 731.165 -0.515 ;
        RECT 729.475 -0.845 729.805 -0.515 ;
        RECT 728.115 -0.845 728.445 -0.515 ;
        RECT 726.755 -0.845 727.085 -0.515 ;
        RECT 725.395 -0.845 725.725 -0.515 ;
        RECT 724.035 -0.845 724.365 -0.515 ;
        RECT 722.675 -0.845 723.005 -0.515 ;
        RECT 721.315 -0.845 721.645 -0.515 ;
        RECT 719.955 -0.845 720.285 -0.515 ;
        RECT 718.595 -0.845 718.925 -0.515 ;
        RECT 717.235 -0.845 717.565 -0.515 ;
        RECT 715.875 -0.845 716.205 -0.515 ;
        RECT 714.515 -0.845 714.845 -0.515 ;
        RECT 713.155 -0.845 713.485 -0.515 ;
        RECT 711.795 -0.845 712.125 -0.515 ;
        RECT 710.435 -0.845 710.765 -0.515 ;
        RECT 709.075 -0.845 709.405 -0.515 ;
        RECT 707.715 -0.845 708.045 -0.515 ;
        RECT 706.355 -0.845 706.685 -0.515 ;
        RECT 704.995 -0.845 705.325 -0.515 ;
        RECT 703.635 -0.845 703.965 -0.515 ;
        RECT 702.275 -0.845 702.605 -0.515 ;
        RECT 700.915 -0.845 701.245 -0.515 ;
        RECT 699.555 -0.845 699.885 -0.515 ;
        RECT 698.195 -0.845 698.525 -0.515 ;
        RECT 696.835 -0.845 697.165 -0.515 ;
        RECT 695.475 -0.845 695.805 -0.515 ;
        RECT 694.115 -0.845 694.445 -0.515 ;
        RECT 692.755 -0.845 693.085 -0.515 ;
        RECT 691.395 -0.845 691.725 -0.515 ;
        RECT 690.035 -0.845 690.365 -0.515 ;
        RECT 688.675 -0.845 689.005 -0.515 ;
        RECT 687.315 -0.845 687.645 -0.515 ;
        RECT 685.955 -0.845 686.285 -0.515 ;
        RECT 684.595 -0.845 684.925 -0.515 ;
        RECT 683.235 -0.845 683.565 -0.515 ;
        RECT 681.875 -0.845 682.205 -0.515 ;
        RECT 680.515 -0.845 680.845 -0.515 ;
        RECT 679.155 -0.845 679.485 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.4 -23.96 226.6 -23.64 ;
        RECT 224.915 -23.965 225.245 -23.635 ;
        RECT 223.555 -23.965 223.885 -23.635 ;
        RECT 222.195 -23.965 222.525 -23.635 ;
        RECT 220.835 -23.965 221.165 -23.635 ;
        RECT 219.475 -23.965 219.805 -23.635 ;
        RECT 216.755 -23.965 217.085 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.08 -28.04 226.6 -27.72 ;
        RECT 224.915 -28.045 225.245 -27.715 ;
        RECT 223.555 -28.045 223.885 -27.715 ;
        RECT 222.195 -28.045 222.525 -27.715 ;
        RECT 220.835 -28.045 221.165 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -34.845 226.605 -34.515 ;
        RECT 219.48 -34.84 226.605 -34.52 ;
        RECT 224.915 -34.845 225.245 -34.515 ;
        RECT 223.555 -34.845 223.885 -34.515 ;
        RECT 222.195 -34.845 222.525 -34.515 ;
        RECT 220.835 -34.845 221.165 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.48 -26.68 230 -26.36 ;
        RECT 228.995 -26.685 229.325 -26.355 ;
        RECT 227.635 -26.685 227.965 -26.355 ;
        RECT 224.915 -26.685 225.245 -26.355 ;
        RECT 223.555 -26.685 223.885 -26.355 ;
        RECT 222.195 -26.685 222.525 -26.355 ;
        RECT 220.835 -26.685 221.165 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.44 -29.4 240.88 -29.08 ;
        RECT 239.875 -29.405 240.205 -29.075 ;
        RECT 238.515 -29.405 238.845 -29.075 ;
        RECT 237.155 -29.405 237.485 -29.075 ;
        RECT 235.795 -29.405 236.125 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.36 -23.96 241.56 -23.64 ;
        RECT 239.875 -23.965 240.205 -23.635 ;
        RECT 238.515 -23.965 238.845 -23.635 ;
        RECT 237.155 -23.965 237.485 -23.635 ;
        RECT 235.795 -23.965 236.125 -23.635 ;
        RECT 234.435 -23.965 234.765 -23.635 ;
        RECT 231.715 -23.965 232.045 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.04 -28.04 241.56 -27.72 ;
        RECT 239.875 -28.045 240.205 -27.715 ;
        RECT 238.515 -28.045 238.845 -27.715 ;
        RECT 237.155 -28.045 237.485 -27.715 ;
        RECT 235.795 -28.045 236.125 -27.715 ;
        RECT 231.715 -28.045 232.045 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 -34.845 241.565 -34.515 ;
        RECT 234.44 -34.84 241.565 -34.52 ;
        RECT 239.875 -34.845 240.205 -34.515 ;
        RECT 238.515 -34.845 238.845 -34.515 ;
        RECT 237.155 -34.845 237.485 -34.515 ;
        RECT 235.795 -34.845 236.125 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.44 -26.68 244.96 -26.36 ;
        RECT 243.955 -26.685 244.285 -26.355 ;
        RECT 242.595 -26.685 242.925 -26.355 ;
        RECT 239.875 -26.685 240.205 -26.355 ;
        RECT 238.515 -26.685 238.845 -26.355 ;
        RECT 237.155 -26.685 237.485 -26.355 ;
        RECT 235.795 -26.685 236.125 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -29.4 255.84 -29.08 ;
        RECT 254.835 -29.405 255.165 -29.075 ;
        RECT 253.475 -29.405 253.805 -29.075 ;
        RECT 252.115 -29.405 252.445 -29.075 ;
        RECT 250.755 -29.405 251.085 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.32 -23.96 256.52 -23.64 ;
        RECT 254.835 -23.965 255.165 -23.635 ;
        RECT 253.475 -23.965 253.805 -23.635 ;
        RECT 252.115 -23.965 252.445 -23.635 ;
        RECT 250.755 -23.965 251.085 -23.635 ;
        RECT 249.395 -23.965 249.725 -23.635 ;
        RECT 246.675 -23.965 247.005 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 246 -28.04 256.52 -27.72 ;
        RECT 254.835 -28.045 255.165 -27.715 ;
        RECT 253.475 -28.045 253.805 -27.715 ;
        RECT 252.115 -28.045 252.445 -27.715 ;
        RECT 250.755 -28.045 251.085 -27.715 ;
        RECT 246.675 -28.045 247.005 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 -34.845 256.525 -34.515 ;
        RECT 249.4 -34.84 256.525 -34.52 ;
        RECT 254.835 -34.845 255.165 -34.515 ;
        RECT 253.475 -34.845 253.805 -34.515 ;
        RECT 252.115 -34.845 252.445 -34.515 ;
        RECT 250.755 -34.845 251.085 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -26.68 259.92 -26.36 ;
        RECT 257.555 -26.685 257.885 -26.355 ;
        RECT 254.835 -26.685 255.165 -26.355 ;
        RECT 253.475 -26.685 253.805 -26.355 ;
        RECT 252.115 -26.685 252.445 -26.355 ;
        RECT 250.755 -26.685 251.085 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.36 -29.4 270.8 -29.08 ;
        RECT 269.795 -29.405 270.125 -29.075 ;
        RECT 268.435 -29.405 268.765 -29.075 ;
        RECT 267.075 -29.405 267.405 -29.075 ;
        RECT 265.715 -29.405 266.045 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 -23.96 271.48 -23.64 ;
        RECT 269.795 -23.965 270.125 -23.635 ;
        RECT 268.435 -23.965 268.765 -23.635 ;
        RECT 267.075 -23.965 267.405 -23.635 ;
        RECT 265.715 -23.965 266.045 -23.635 ;
        RECT 264.355 -23.965 264.685 -23.635 ;
        RECT 261.635 -23.965 261.965 -23.635 ;
        RECT 260.275 -23.965 260.605 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.28 -28.04 271.48 -27.72 ;
        RECT 269.795 -28.045 270.125 -27.715 ;
        RECT 268.435 -28.045 268.765 -27.715 ;
        RECT 267.075 -28.045 267.405 -27.715 ;
        RECT 265.715 -28.045 266.045 -27.715 ;
        RECT 261.635 -28.045 261.965 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 -34.845 271.485 -34.515 ;
        RECT 264.36 -34.84 271.485 -34.52 ;
        RECT 269.795 -34.845 270.125 -34.515 ;
        RECT 268.435 -34.845 268.765 -34.515 ;
        RECT 267.075 -34.845 267.405 -34.515 ;
        RECT 265.715 -34.845 266.045 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.36 -26.68 274.88 -26.36 ;
        RECT 272.515 -26.685 272.845 -26.355 ;
        RECT 269.795 -26.685 270.125 -26.355 ;
        RECT 268.435 -26.685 268.765 -26.355 ;
        RECT 267.075 -26.685 267.405 -26.355 ;
        RECT 265.715 -26.685 266.045 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.32 -29.4 285.76 -29.08 ;
        RECT 284.755 -29.405 285.085 -29.075 ;
        RECT 283.395 -29.405 283.725 -29.075 ;
        RECT 282.035 -29.405 282.365 -29.075 ;
        RECT 280.675 -29.405 281.005 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.56 -23.96 286.44 -23.64 ;
        RECT 284.755 -23.965 285.085 -23.635 ;
        RECT 283.395 -23.965 283.725 -23.635 ;
        RECT 282.035 -23.965 282.365 -23.635 ;
        RECT 280.675 -23.965 281.005 -23.635 ;
        RECT 279.315 -23.965 279.645 -23.635 ;
        RECT 276.595 -23.965 276.925 -23.635 ;
        RECT 275.235 -23.965 275.565 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.24 -28.04 286.44 -27.72 ;
        RECT 284.755 -28.045 285.085 -27.715 ;
        RECT 283.395 -28.045 283.725 -27.715 ;
        RECT 282.035 -28.045 282.365 -27.715 ;
        RECT 280.675 -28.045 281.005 -27.715 ;
        RECT 276.595 -28.045 276.925 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 -34.845 286.445 -34.515 ;
        RECT 279.32 -34.84 286.445 -34.52 ;
        RECT 284.755 -34.845 285.085 -34.515 ;
        RECT 283.395 -34.845 283.725 -34.515 ;
        RECT 282.035 -34.845 282.365 -34.515 ;
        RECT 280.675 -34.845 281.005 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.32 -26.68 289.84 -26.36 ;
        RECT 287.475 -26.685 287.805 -26.355 ;
        RECT 284.755 -26.685 285.085 -26.355 ;
        RECT 283.395 -26.685 283.725 -26.355 ;
        RECT 282.035 -26.685 282.365 -26.355 ;
        RECT 280.675 -26.685 281.005 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.52 -23.96 300.72 -23.64 ;
        RECT 298.355 -23.965 298.685 -23.635 ;
        RECT 296.995 -23.965 297.325 -23.635 ;
        RECT 295.635 -23.965 295.965 -23.635 ;
        RECT 294.275 -23.965 294.605 -23.635 ;
        RECT 291.555 -23.965 291.885 -23.635 ;
        RECT 290.195 -23.965 290.525 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -28.04 300.72 -27.72 ;
        RECT 298.355 -28.045 298.685 -27.715 ;
        RECT 296.995 -28.045 297.325 -27.715 ;
        RECT 295.635 -28.045 295.965 -27.715 ;
        RECT 291.555 -28.045 291.885 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.28 -29.4 300.72 -29.08 ;
        RECT 298.355 -29.405 298.685 -29.075 ;
        RECT 296.995 -29.405 297.325 -29.075 ;
        RECT 295.635 -29.405 295.965 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.28 -34.84 300.72 -34.52 ;
        RECT 299.715 -34.845 300.045 -34.515 ;
        RECT 298.355 -34.845 298.685 -34.515 ;
        RECT 296.995 -34.845 297.325 -34.515 ;
        RECT 295.635 -34.845 295.965 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.28 -26.68 304.8 -26.36 ;
        RECT 302.435 -26.685 302.765 -26.355 ;
        RECT 298.355 -26.685 298.685 -26.355 ;
        RECT 296.995 -26.685 297.325 -26.355 ;
        RECT 295.635 -26.685 295.965 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.24 -29.4 315 -29.08 ;
        RECT 313.315 -29.405 313.645 -29.075 ;
        RECT 311.955 -29.405 312.285 -29.075 ;
        RECT 310.595 -29.405 310.925 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.48 -23.96 315.68 -23.64 ;
        RECT 313.315 -23.965 313.645 -23.635 ;
        RECT 311.955 -23.965 312.285 -23.635 ;
        RECT 310.595 -23.965 310.925 -23.635 ;
        RECT 309.235 -23.965 309.565 -23.635 ;
        RECT 306.515 -23.965 306.845 -23.635 ;
        RECT 305.155 -23.965 305.485 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.16 -28.04 315.68 -27.72 ;
        RECT 313.315 -28.045 313.645 -27.715 ;
        RECT 311.955 -28.045 312.285 -27.715 ;
        RECT 310.595 -28.045 310.925 -27.715 ;
        RECT 306.515 -28.045 306.845 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.24 -34.84 315.68 -34.52 ;
        RECT 314.675 -34.845 315.005 -34.515 ;
        RECT 313.315 -34.845 313.645 -34.515 ;
        RECT 311.955 -34.845 312.285 -34.515 ;
        RECT 310.595 -34.845 310.925 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.24 -26.68 319.76 -26.36 ;
        RECT 317.395 -26.685 317.725 -26.355 ;
        RECT 313.315 -26.685 313.645 -26.355 ;
        RECT 311.955 -26.685 312.285 -26.355 ;
        RECT 310.595 -26.685 310.925 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.2 -29.4 329.96 -29.08 ;
        RECT 328.275 -29.405 328.605 -29.075 ;
        RECT 326.915 -29.405 327.245 -29.075 ;
        RECT 325.555 -29.405 325.885 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.44 -23.96 330.64 -23.64 ;
        RECT 328.275 -23.965 328.605 -23.635 ;
        RECT 326.915 -23.965 327.245 -23.635 ;
        RECT 325.555 -23.965 325.885 -23.635 ;
        RECT 324.195 -23.965 324.525 -23.635 ;
        RECT 321.475 -23.965 321.805 -23.635 ;
        RECT 320.115 -23.965 320.445 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.12 -28.04 330.64 -27.72 ;
        RECT 328.275 -28.045 328.605 -27.715 ;
        RECT 326.915 -28.045 327.245 -27.715 ;
        RECT 325.555 -28.045 325.885 -27.715 ;
        RECT 321.475 -28.045 321.805 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.2 -34.84 330.64 -34.52 ;
        RECT 329.635 -34.845 329.965 -34.515 ;
        RECT 328.275 -34.845 328.605 -34.515 ;
        RECT 326.915 -34.845 327.245 -34.515 ;
        RECT 325.555 -34.845 325.885 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.2 -26.68 334.72 -26.36 ;
        RECT 332.355 -26.685 332.685 -26.355 ;
        RECT 328.275 -26.685 328.605 -26.355 ;
        RECT 326.915 -26.685 327.245 -26.355 ;
        RECT 325.555 -26.685 325.885 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -29.4 344.92 -29.08 ;
        RECT 343.235 -29.405 343.565 -29.075 ;
        RECT 341.875 -29.405 342.205 -29.075 ;
        RECT 340.515 -29.405 340.845 -29.075 ;
        RECT 339.155 -29.405 339.485 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.4 -23.96 345.6 -23.64 ;
        RECT 343.235 -23.965 343.565 -23.635 ;
        RECT 341.875 -23.965 342.205 -23.635 ;
        RECT 340.515 -23.965 340.845 -23.635 ;
        RECT 339.155 -23.965 339.485 -23.635 ;
        RECT 336.435 -23.965 336.765 -23.635 ;
        RECT 335.075 -23.965 335.405 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.08 -28.04 345.6 -27.72 ;
        RECT 343.235 -28.045 343.565 -27.715 ;
        RECT 341.875 -28.045 342.205 -27.715 ;
        RECT 340.515 -28.045 340.845 -27.715 ;
        RECT 339.155 -28.045 339.485 -27.715 ;
        RECT 336.435 -28.045 336.765 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -34.84 345.6 -34.52 ;
        RECT 344.595 -34.845 344.925 -34.515 ;
        RECT 343.235 -34.845 343.565 -34.515 ;
        RECT 341.875 -34.845 342.205 -34.515 ;
        RECT 340.515 -34.845 340.845 -34.515 ;
        RECT 339.155 -34.845 339.485 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -26.68 349.68 -26.36 ;
        RECT 347.315 -26.685 347.645 -26.355 ;
        RECT 343.235 -26.685 343.565 -26.355 ;
        RECT 341.875 -26.685 342.205 -26.355 ;
        RECT 340.515 -26.685 340.845 -26.355 ;
        RECT 339.155 -26.685 339.485 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.44 -29.4 359.88 -29.08 ;
        RECT 358.195 -29.405 358.525 -29.075 ;
        RECT 356.835 -29.405 357.165 -29.075 ;
        RECT 355.475 -29.405 355.805 -29.075 ;
        RECT 354.115 -29.405 354.445 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.36 -23.96 360.56 -23.64 ;
        RECT 358.195 -23.965 358.525 -23.635 ;
        RECT 356.835 -23.965 357.165 -23.635 ;
        RECT 355.475 -23.965 355.805 -23.635 ;
        RECT 354.115 -23.965 354.445 -23.635 ;
        RECT 351.395 -23.965 351.725 -23.635 ;
        RECT 350.035 -23.965 350.365 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.04 -28.04 360.56 -27.72 ;
        RECT 358.195 -28.045 358.525 -27.715 ;
        RECT 356.835 -28.045 357.165 -27.715 ;
        RECT 355.475 -28.045 355.805 -27.715 ;
        RECT 354.115 -28.045 354.445 -27.715 ;
        RECT 351.395 -28.045 351.725 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.44 -34.84 360.56 -34.52 ;
        RECT 359.555 -34.845 359.885 -34.515 ;
        RECT 358.195 -34.845 358.525 -34.515 ;
        RECT 356.835 -34.845 357.165 -34.515 ;
        RECT 355.475 -34.845 355.805 -34.515 ;
        RECT 354.115 -34.845 354.445 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.44 -26.68 364.64 -26.36 ;
        RECT 362.275 -26.685 362.605 -26.355 ;
        RECT 358.195 -26.685 358.525 -26.355 ;
        RECT 356.835 -26.685 357.165 -26.355 ;
        RECT 355.475 -26.685 355.805 -26.355 ;
        RECT 354.115 -26.685 354.445 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.4 -29.4 374.84 -29.08 ;
        RECT 373.155 -29.405 373.485 -29.075 ;
        RECT 371.795 -29.405 372.125 -29.075 ;
        RECT 370.435 -29.405 370.765 -29.075 ;
        RECT 369.075 -29.405 369.405 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.32 -23.96 375.52 -23.64 ;
        RECT 373.155 -23.965 373.485 -23.635 ;
        RECT 371.795 -23.965 372.125 -23.635 ;
        RECT 370.435 -23.965 370.765 -23.635 ;
        RECT 369.075 -23.965 369.405 -23.635 ;
        RECT 364.995 -23.965 365.325 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 365 -28.04 375.52 -27.72 ;
        RECT 373.155 -28.045 373.485 -27.715 ;
        RECT 371.795 -28.045 372.125 -27.715 ;
        RECT 370.435 -28.045 370.765 -27.715 ;
        RECT 369.075 -28.045 369.405 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.4 -34.84 375.52 -34.52 ;
        RECT 374.515 -34.845 374.845 -34.515 ;
        RECT 373.155 -34.845 373.485 -34.515 ;
        RECT 371.795 -34.845 372.125 -34.515 ;
        RECT 370.435 -34.845 370.765 -34.515 ;
        RECT 369.075 -34.845 369.405 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.4 -26.68 379.6 -26.36 ;
        RECT 377.235 -26.685 377.565 -26.355 ;
        RECT 373.155 -26.685 373.485 -26.355 ;
        RECT 371.795 -26.685 372.125 -26.355 ;
        RECT 370.435 -26.685 370.765 -26.355 ;
        RECT 369.075 -26.685 369.405 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.36 -29.4 389.8 -29.08 ;
        RECT 388.115 -29.405 388.445 -29.075 ;
        RECT 386.755 -29.405 387.085 -29.075 ;
        RECT 385.395 -29.405 385.725 -29.075 ;
        RECT 384.035 -29.405 384.365 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.28 -23.96 390.48 -23.64 ;
        RECT 388.115 -23.965 388.445 -23.635 ;
        RECT 386.755 -23.965 387.085 -23.635 ;
        RECT 385.395 -23.965 385.725 -23.635 ;
        RECT 384.035 -23.965 384.365 -23.635 ;
        RECT 379.955 -23.965 380.285 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.96 -28.04 390.48 -27.72 ;
        RECT 388.115 -28.045 388.445 -27.715 ;
        RECT 386.755 -28.045 387.085 -27.715 ;
        RECT 385.395 -28.045 385.725 -27.715 ;
        RECT 384.035 -28.045 384.365 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.36 -34.84 390.48 -34.52 ;
        RECT 389.475 -34.845 389.805 -34.515 ;
        RECT 388.115 -34.845 388.445 -34.515 ;
        RECT 386.755 -34.845 387.085 -34.515 ;
        RECT 385.395 -34.845 385.725 -34.515 ;
        RECT 384.035 -34.845 384.365 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.36 -26.68 393.88 -26.36 ;
        RECT 392.195 -26.685 392.525 -26.355 ;
        RECT 388.115 -26.685 388.445 -26.355 ;
        RECT 386.755 -26.685 387.085 -26.355 ;
        RECT 385.395 -26.685 385.725 -26.355 ;
        RECT 384.035 -26.685 384.365 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.32 -29.4 404.76 -29.08 ;
        RECT 403.075 -29.405 403.405 -29.075 ;
        RECT 401.715 -29.405 402.045 -29.075 ;
        RECT 400.355 -29.405 400.685 -29.075 ;
        RECT 398.995 -29.405 399.325 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.24 -23.96 405.44 -23.64 ;
        RECT 403.075 -23.965 403.405 -23.635 ;
        RECT 401.715 -23.965 402.045 -23.635 ;
        RECT 400.355 -23.965 400.685 -23.635 ;
        RECT 398.995 -23.965 399.325 -23.635 ;
        RECT 394.915 -23.965 395.245 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.92 -28.04 405.44 -27.72 ;
        RECT 403.075 -28.045 403.405 -27.715 ;
        RECT 401.715 -28.045 402.045 -27.715 ;
        RECT 400.355 -28.045 400.685 -27.715 ;
        RECT 398.995 -28.045 399.325 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.32 -34.84 405.44 -34.52 ;
        RECT 404.435 -34.845 404.765 -34.515 ;
        RECT 403.075 -34.845 403.405 -34.515 ;
        RECT 401.715 -34.845 402.045 -34.515 ;
        RECT 400.355 -34.845 400.685 -34.515 ;
        RECT 398.995 -34.845 399.325 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.32 -26.68 408.84 -26.36 ;
        RECT 407.155 -26.685 407.485 -26.355 ;
        RECT 403.075 -26.685 403.405 -26.355 ;
        RECT 401.715 -26.685 402.045 -26.355 ;
        RECT 400.355 -26.685 400.685 -26.355 ;
        RECT 398.995 -26.685 399.325 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.28 -29.4 419.72 -29.08 ;
        RECT 418.035 -29.405 418.365 -29.075 ;
        RECT 416.675 -29.405 417.005 -29.075 ;
        RECT 415.315 -29.405 415.645 -29.075 ;
        RECT 413.955 -29.405 414.285 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.2 -23.96 420.4 -23.64 ;
        RECT 418.035 -23.965 418.365 -23.635 ;
        RECT 416.675 -23.965 417.005 -23.635 ;
        RECT 415.315 -23.965 415.645 -23.635 ;
        RECT 413.955 -23.965 414.285 -23.635 ;
        RECT 409.875 -23.965 410.205 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.88 -28.04 420.4 -27.72 ;
        RECT 418.035 -28.045 418.365 -27.715 ;
        RECT 416.675 -28.045 417.005 -27.715 ;
        RECT 415.315 -28.045 415.645 -27.715 ;
        RECT 413.955 -28.045 414.285 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.28 -34.84 420.4 -34.52 ;
        RECT 419.395 -34.845 419.725 -34.515 ;
        RECT 418.035 -34.845 418.365 -34.515 ;
        RECT 416.675 -34.845 417.005 -34.515 ;
        RECT 415.315 -34.845 415.645 -34.515 ;
        RECT 413.955 -34.845 414.285 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.28 -26.68 423.8 -26.36 ;
        RECT 422.115 -26.685 422.445 -26.355 ;
        RECT 418.035 -26.685 418.365 -26.355 ;
        RECT 416.675 -26.685 417.005 -26.355 ;
        RECT 415.315 -26.685 415.645 -26.355 ;
        RECT 413.955 -26.685 414.285 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.24 -29.4 434.68 -29.08 ;
        RECT 432.995 -29.405 433.325 -29.075 ;
        RECT 431.635 -29.405 431.965 -29.075 ;
        RECT 430.275 -29.405 430.605 -29.075 ;
        RECT 428.915 -29.405 429.245 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.16 -23.96 435.36 -23.64 ;
        RECT 432.995 -23.965 433.325 -23.635 ;
        RECT 431.635 -23.965 431.965 -23.635 ;
        RECT 430.275 -23.965 430.605 -23.635 ;
        RECT 428.915 -23.965 429.245 -23.635 ;
        RECT 424.835 -23.965 425.165 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.16 -28.04 435.36 -27.72 ;
        RECT 432.995 -28.045 433.325 -27.715 ;
        RECT 431.635 -28.045 431.965 -27.715 ;
        RECT 430.275 -28.045 430.605 -27.715 ;
        RECT 428.915 -28.045 429.245 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.24 -34.84 435.36 -34.52 ;
        RECT 434.355 -34.845 434.685 -34.515 ;
        RECT 432.995 -34.845 433.325 -34.515 ;
        RECT 431.635 -34.845 431.965 -34.515 ;
        RECT 430.275 -34.845 430.605 -34.515 ;
        RECT 428.915 -34.845 429.245 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.24 -26.68 438.76 -26.36 ;
        RECT 437.075 -26.685 437.405 -26.355 ;
        RECT 432.995 -26.685 433.325 -26.355 ;
        RECT 431.635 -26.685 431.965 -26.355 ;
        RECT 430.275 -26.685 430.605 -26.355 ;
        RECT 428.915 -26.685 429.245 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.2 -29.4 449.64 -29.08 ;
        RECT 447.955 -29.405 448.285 -29.075 ;
        RECT 446.595 -29.405 446.925 -29.075 ;
        RECT 445.235 -29.405 445.565 -29.075 ;
        RECT 443.875 -29.405 444.205 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.44 -23.96 450.32 -23.64 ;
        RECT 447.955 -23.965 448.285 -23.635 ;
        RECT 446.595 -23.965 446.925 -23.635 ;
        RECT 445.235 -23.965 445.565 -23.635 ;
        RECT 443.875 -23.965 444.205 -23.635 ;
        RECT 439.795 -23.965 440.125 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.12 -28.04 450.32 -27.72 ;
        RECT 447.955 -28.045 448.285 -27.715 ;
        RECT 446.595 -28.045 446.925 -27.715 ;
        RECT 445.235 -28.045 445.565 -27.715 ;
        RECT 443.875 -28.045 444.205 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.2 -34.84 450.32 -34.52 ;
        RECT 449.315 -34.845 449.645 -34.515 ;
        RECT 447.955 -34.845 448.285 -34.515 ;
        RECT 446.595 -34.845 446.925 -34.515 ;
        RECT 445.235 -34.845 445.565 -34.515 ;
        RECT 443.875 -34.845 444.205 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.2 -26.68 453.72 -26.36 ;
        RECT 452.035 -26.685 452.365 -26.355 ;
        RECT 447.955 -26.685 448.285 -26.355 ;
        RECT 446.595 -26.685 446.925 -26.355 ;
        RECT 445.235 -26.685 445.565 -26.355 ;
        RECT 443.875 -26.685 444.205 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -23.96 464.6 -23.64 ;
        RECT 462.915 -23.965 463.245 -23.635 ;
        RECT 461.555 -23.965 461.885 -23.635 ;
        RECT 460.195 -23.965 460.525 -23.635 ;
        RECT 458.835 -23.965 459.165 -23.635 ;
        RECT 454.755 -23.965 455.085 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.08 -28.04 464.6 -27.72 ;
        RECT 462.915 -28.045 463.245 -27.715 ;
        RECT 461.555 -28.045 461.885 -27.715 ;
        RECT 460.195 -28.045 460.525 -27.715 ;
        RECT 458.835 -28.045 459.165 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.16 -29.4 464.6 -29.08 ;
        RECT 462.915 -29.405 463.245 -29.075 ;
        RECT 461.555 -29.405 461.885 -29.075 ;
        RECT 460.195 -29.405 460.525 -29.075 ;
        RECT 458.835 -29.405 459.165 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 464.275 -34.845 464.605 -34.515 ;
        RECT 458.16 -34.84 464.605 -34.52 ;
        RECT 462.915 -34.845 463.245 -34.515 ;
        RECT 461.555 -34.845 461.885 -34.515 ;
        RECT 460.195 -34.845 460.525 -34.515 ;
        RECT 458.835 -34.845 459.165 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.16 -26.68 468.68 -26.36 ;
        RECT 466.995 -26.685 467.325 -26.355 ;
        RECT 462.915 -26.685 463.245 -26.355 ;
        RECT 461.555 -26.685 461.885 -26.355 ;
        RECT 460.195 -26.685 460.525 -26.355 ;
        RECT 458.835 -26.685 459.165 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.12 -29.4 478.88 -29.08 ;
        RECT 477.875 -29.405 478.205 -29.075 ;
        RECT 476.515 -29.405 476.845 -29.075 ;
        RECT 475.155 -29.405 475.485 -29.075 ;
        RECT 473.795 -29.405 474.125 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.36 -23.96 479.56 -23.64 ;
        RECT 477.875 -23.965 478.205 -23.635 ;
        RECT 476.515 -23.965 476.845 -23.635 ;
        RECT 475.155 -23.965 475.485 -23.635 ;
        RECT 473.795 -23.965 474.125 -23.635 ;
        RECT 469.715 -23.965 470.045 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.04 -28.04 479.56 -27.72 ;
        RECT 477.875 -28.045 478.205 -27.715 ;
        RECT 476.515 -28.045 476.845 -27.715 ;
        RECT 475.155 -28.045 475.485 -27.715 ;
        RECT 473.795 -28.045 474.125 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 479.235 -34.845 479.565 -34.515 ;
        RECT 473.12 -34.84 479.565 -34.52 ;
        RECT 477.875 -34.845 478.205 -34.515 ;
        RECT 476.515 -34.845 476.845 -34.515 ;
        RECT 475.155 -34.845 475.485 -34.515 ;
        RECT 473.795 -34.845 474.125 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.12 -26.68 483.64 -26.36 ;
        RECT 481.955 -26.685 482.285 -26.355 ;
        RECT 480.595 -26.685 480.925 -26.355 ;
        RECT 477.875 -26.685 478.205 -26.355 ;
        RECT 476.515 -26.685 476.845 -26.355 ;
        RECT 475.155 -26.685 475.485 -26.355 ;
        RECT 473.795 -26.685 474.125 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.08 -29.4 493.84 -29.08 ;
        RECT 492.835 -29.405 493.165 -29.075 ;
        RECT 491.475 -29.405 491.805 -29.075 ;
        RECT 490.115 -29.405 490.445 -29.075 ;
        RECT 488.755 -29.405 489.085 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.32 -23.96 494.52 -23.64 ;
        RECT 492.835 -23.965 493.165 -23.635 ;
        RECT 491.475 -23.965 491.805 -23.635 ;
        RECT 490.115 -23.965 490.445 -23.635 ;
        RECT 488.755 -23.965 489.085 -23.635 ;
        RECT 484.675 -23.965 485.005 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 484 -28.04 494.52 -27.72 ;
        RECT 492.835 -28.045 493.165 -27.715 ;
        RECT 491.475 -28.045 491.805 -27.715 ;
        RECT 490.115 -28.045 490.445 -27.715 ;
        RECT 488.755 -28.045 489.085 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 494.195 -34.845 494.525 -34.515 ;
        RECT 488.08 -34.84 494.525 -34.52 ;
        RECT 492.835 -34.845 493.165 -34.515 ;
        RECT 491.475 -34.845 491.805 -34.515 ;
        RECT 490.115 -34.845 490.445 -34.515 ;
        RECT 488.755 -34.845 489.085 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.08 -26.68 498.6 -26.36 ;
        RECT 496.915 -26.685 497.245 -26.355 ;
        RECT 495.555 -26.685 495.885 -26.355 ;
        RECT 492.835 -26.685 493.165 -26.355 ;
        RECT 491.475 -26.685 491.805 -26.355 ;
        RECT 490.115 -26.685 490.445 -26.355 ;
        RECT 488.755 -26.685 489.085 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.04 -29.4 508.8 -29.08 ;
        RECT 507.795 -29.405 508.125 -29.075 ;
        RECT 506.435 -29.405 506.765 -29.075 ;
        RECT 505.075 -29.405 505.405 -29.075 ;
        RECT 503.715 -29.405 504.045 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.28 -23.96 509.48 -23.64 ;
        RECT 507.795 -23.965 508.125 -23.635 ;
        RECT 506.435 -23.965 506.765 -23.635 ;
        RECT 505.075 -23.965 505.405 -23.635 ;
        RECT 503.715 -23.965 504.045 -23.635 ;
        RECT 499.635 -23.965 499.965 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.96 -28.04 509.48 -27.72 ;
        RECT 507.795 -28.045 508.125 -27.715 ;
        RECT 506.435 -28.045 506.765 -27.715 ;
        RECT 505.075 -28.045 505.405 -27.715 ;
        RECT 503.715 -28.045 504.045 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 509.155 -34.845 509.485 -34.515 ;
        RECT 503.04 -34.84 509.485 -34.52 ;
        RECT 507.795 -34.845 508.125 -34.515 ;
        RECT 506.435 -34.845 506.765 -34.515 ;
        RECT 505.075 -34.845 505.405 -34.515 ;
        RECT 503.715 -34.845 504.045 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.04 -26.68 513.56 -26.36 ;
        RECT 511.875 -26.685 512.205 -26.355 ;
        RECT 510.515 -26.685 510.845 -26.355 ;
        RECT 507.795 -26.685 508.125 -26.355 ;
        RECT 506.435 -26.685 506.765 -26.355 ;
        RECT 505.075 -26.685 505.405 -26.355 ;
        RECT 503.715 -26.685 504.045 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 518 -29.4 523.76 -29.08 ;
        RECT 522.755 -29.405 523.085 -29.075 ;
        RECT 521.395 -29.405 521.725 -29.075 ;
        RECT 520.035 -29.405 520.365 -29.075 ;
        RECT 518.675 -29.405 519.005 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.24 -23.96 524.44 -23.64 ;
        RECT 522.755 -23.965 523.085 -23.635 ;
        RECT 521.395 -23.965 521.725 -23.635 ;
        RECT 520.035 -23.965 520.365 -23.635 ;
        RECT 518.675 -23.965 519.005 -23.635 ;
        RECT 517.315 -23.965 517.645 -23.635 ;
        RECT 514.595 -23.965 514.925 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.92 -28.04 524.44 -27.72 ;
        RECT 522.755 -28.045 523.085 -27.715 ;
        RECT 521.395 -28.045 521.725 -27.715 ;
        RECT 520.035 -28.045 520.365 -27.715 ;
        RECT 518.675 -28.045 519.005 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 524.115 -34.845 524.445 -34.515 ;
        RECT 518 -34.84 524.445 -34.52 ;
        RECT 522.755 -34.845 523.085 -34.515 ;
        RECT 521.395 -34.845 521.725 -34.515 ;
        RECT 520.035 -34.845 520.365 -34.515 ;
        RECT 518.675 -34.845 519.005 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 518 -26.68 528.52 -26.36 ;
        RECT 526.835 -26.685 527.165 -26.355 ;
        RECT 525.475 -26.685 525.805 -26.355 ;
        RECT 522.755 -26.685 523.085 -26.355 ;
        RECT 521.395 -26.685 521.725 -26.355 ;
        RECT 520.035 -26.685 520.365 -26.355 ;
        RECT 518.675 -26.685 519.005 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.28 -29.4 538.72 -29.08 ;
        RECT 537.715 -29.405 538.045 -29.075 ;
        RECT 536.355 -29.405 536.685 -29.075 ;
        RECT 534.995 -29.405 535.325 -29.075 ;
        RECT 533.635 -29.405 533.965 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.2 -23.96 539.4 -23.64 ;
        RECT 537.715 -23.965 538.045 -23.635 ;
        RECT 536.355 -23.965 536.685 -23.635 ;
        RECT 534.995 -23.965 535.325 -23.635 ;
        RECT 533.635 -23.965 533.965 -23.635 ;
        RECT 532.275 -23.965 532.605 -23.635 ;
        RECT 529.555 -23.965 529.885 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.88 -28.04 539.4 -27.72 ;
        RECT 537.715 -28.045 538.045 -27.715 ;
        RECT 536.355 -28.045 536.685 -27.715 ;
        RECT 534.995 -28.045 535.325 -27.715 ;
        RECT 533.635 -28.045 533.965 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 539.075 -34.845 539.405 -34.515 ;
        RECT 532.28 -34.84 539.405 -34.52 ;
        RECT 537.715 -34.845 538.045 -34.515 ;
        RECT 536.355 -34.845 536.685 -34.515 ;
        RECT 534.995 -34.845 535.325 -34.515 ;
        RECT 533.635 -34.845 533.965 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.28 -26.68 543.48 -26.36 ;
        RECT 541.795 -26.685 542.125 -26.355 ;
        RECT 540.435 -26.685 540.765 -26.355 ;
        RECT 537.715 -26.685 538.045 -26.355 ;
        RECT 536.355 -26.685 536.685 -26.355 ;
        RECT 534.995 -26.685 535.325 -26.355 ;
        RECT 533.635 -26.685 533.965 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.24 -29.4 553.68 -29.08 ;
        RECT 552.675 -29.405 553.005 -29.075 ;
        RECT 551.315 -29.405 551.645 -29.075 ;
        RECT 549.955 -29.405 550.285 -29.075 ;
        RECT 548.595 -29.405 548.925 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.16 -23.96 554.36 -23.64 ;
        RECT 552.675 -23.965 553.005 -23.635 ;
        RECT 551.315 -23.965 551.645 -23.635 ;
        RECT 549.955 -23.965 550.285 -23.635 ;
        RECT 548.595 -23.965 548.925 -23.635 ;
        RECT 547.235 -23.965 547.565 -23.635 ;
        RECT 544.515 -23.965 544.845 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.84 -28.04 554.36 -27.72 ;
        RECT 552.675 -28.045 553.005 -27.715 ;
        RECT 551.315 -28.045 551.645 -27.715 ;
        RECT 549.955 -28.045 550.285 -27.715 ;
        RECT 548.595 -28.045 548.925 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 554.035 -34.845 554.365 -34.515 ;
        RECT 547.24 -34.84 554.365 -34.52 ;
        RECT 552.675 -34.845 553.005 -34.515 ;
        RECT 551.315 -34.845 551.645 -34.515 ;
        RECT 549.955 -34.845 550.285 -34.515 ;
        RECT 548.595 -34.845 548.925 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.24 -26.68 558.44 -26.36 ;
        RECT 556.755 -26.685 557.085 -26.355 ;
        RECT 555.395 -26.685 555.725 -26.355 ;
        RECT 552.675 -26.685 553.005 -26.355 ;
        RECT 551.315 -26.685 551.645 -26.355 ;
        RECT 549.955 -26.685 550.285 -26.355 ;
        RECT 548.595 -26.685 548.925 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -29.4 568.64 -29.08 ;
        RECT 567.635 -29.405 567.965 -29.075 ;
        RECT 566.275 -29.405 566.605 -29.075 ;
        RECT 564.915 -29.405 565.245 -29.075 ;
        RECT 563.555 -29.405 563.885 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.12 -23.96 569.32 -23.64 ;
        RECT 567.635 -23.965 567.965 -23.635 ;
        RECT 566.275 -23.965 566.605 -23.635 ;
        RECT 564.915 -23.965 565.245 -23.635 ;
        RECT 563.555 -23.965 563.885 -23.635 ;
        RECT 562.195 -23.965 562.525 -23.635 ;
        RECT 559.475 -23.965 559.805 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.8 -28.04 569.32 -27.72 ;
        RECT 567.635 -28.045 567.965 -27.715 ;
        RECT 566.275 -28.045 566.605 -27.715 ;
        RECT 564.915 -28.045 565.245 -27.715 ;
        RECT 563.555 -28.045 563.885 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 568.995 -34.845 569.325 -34.515 ;
        RECT 562.2 -34.84 569.325 -34.52 ;
        RECT 567.635 -34.845 567.965 -34.515 ;
        RECT 566.275 -34.845 566.605 -34.515 ;
        RECT 564.915 -34.845 565.245 -34.515 ;
        RECT 563.555 -34.845 563.885 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -26.68 572.72 -26.36 ;
        RECT 571.715 -26.685 572.045 -26.355 ;
        RECT 570.355 -26.685 570.685 -26.355 ;
        RECT 567.635 -26.685 567.965 -26.355 ;
        RECT 566.275 -26.685 566.605 -26.355 ;
        RECT 564.915 -26.685 565.245 -26.355 ;
        RECT 563.555 -26.685 563.885 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.16 -29.4 583.6 -29.08 ;
        RECT 582.595 -29.405 582.925 -29.075 ;
        RECT 581.235 -29.405 581.565 -29.075 ;
        RECT 579.875 -29.405 580.205 -29.075 ;
        RECT 578.515 -29.405 578.845 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.08 -23.96 584.28 -23.64 ;
        RECT 582.595 -23.965 582.925 -23.635 ;
        RECT 581.235 -23.965 581.565 -23.635 ;
        RECT 579.875 -23.965 580.205 -23.635 ;
        RECT 578.515 -23.965 578.845 -23.635 ;
        RECT 577.155 -23.965 577.485 -23.635 ;
        RECT 574.435 -23.965 574.765 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.76 -28.04 584.28 -27.72 ;
        RECT 582.595 -28.045 582.925 -27.715 ;
        RECT 581.235 -28.045 581.565 -27.715 ;
        RECT 579.875 -28.045 580.205 -27.715 ;
        RECT 578.515 -28.045 578.845 -27.715 ;
        RECT 574.435 -28.045 574.765 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 583.955 -34.845 584.285 -34.515 ;
        RECT 577.16 -34.84 584.285 -34.52 ;
        RECT 582.595 -34.845 582.925 -34.515 ;
        RECT 581.235 -34.845 581.565 -34.515 ;
        RECT 579.875 -34.845 580.205 -34.515 ;
        RECT 578.515 -34.845 578.845 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.16 -26.68 587.68 -26.36 ;
        RECT 586.675 -26.685 587.005 -26.355 ;
        RECT 585.315 -26.685 585.645 -26.355 ;
        RECT 582.595 -26.685 582.925 -26.355 ;
        RECT 581.235 -26.685 581.565 -26.355 ;
        RECT 579.875 -26.685 580.205 -26.355 ;
        RECT 578.515 -26.685 578.845 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.12 -29.4 598.56 -29.08 ;
        RECT 597.555 -29.405 597.885 -29.075 ;
        RECT 596.195 -29.405 596.525 -29.075 ;
        RECT 594.835 -29.405 595.165 -29.075 ;
        RECT 593.475 -29.405 593.805 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.035 -23.96 599.24 -23.64 ;
        RECT 597.555 -23.965 597.885 -23.635 ;
        RECT 596.195 -23.965 596.525 -23.635 ;
        RECT 594.835 -23.965 595.165 -23.635 ;
        RECT 593.475 -23.965 593.805 -23.635 ;
        RECT 592.115 -23.965 592.445 -23.635 ;
        RECT 589.395 -23.965 589.725 -23.635 ;
        RECT 588.035 -23.965 588.365 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.72 -28.04 599.24 -27.72 ;
        RECT 597.555 -28.045 597.885 -27.715 ;
        RECT 596.195 -28.045 596.525 -27.715 ;
        RECT 594.835 -28.045 595.165 -27.715 ;
        RECT 593.475 -28.045 593.805 -27.715 ;
        RECT 589.395 -28.045 589.725 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 598.915 -34.845 599.245 -34.515 ;
        RECT 592.12 -34.84 599.245 -34.52 ;
        RECT 597.555 -34.845 597.885 -34.515 ;
        RECT 596.195 -34.845 596.525 -34.515 ;
        RECT 594.835 -34.845 595.165 -34.515 ;
        RECT 593.475 -34.845 593.805 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.12 -26.68 602.64 -26.36 ;
        RECT 600.275 -26.685 600.605 -26.355 ;
        RECT 597.555 -26.685 597.885 -26.355 ;
        RECT 596.195 -26.685 596.525 -26.355 ;
        RECT 594.835 -26.685 595.165 -26.355 ;
        RECT 593.475 -26.685 593.805 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.08 -29.4 613.52 -29.08 ;
        RECT 612.515 -29.405 612.845 -29.075 ;
        RECT 611.155 -29.405 611.485 -29.075 ;
        RECT 609.795 -29.405 610.125 -29.075 ;
        RECT 608.435 -29.405 608.765 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.32 -23.96 614.2 -23.64 ;
        RECT 612.515 -23.965 612.845 -23.635 ;
        RECT 611.155 -23.965 611.485 -23.635 ;
        RECT 609.795 -23.965 610.125 -23.635 ;
        RECT 608.435 -23.965 608.765 -23.635 ;
        RECT 607.075 -23.965 607.405 -23.635 ;
        RECT 604.355 -23.965 604.685 -23.635 ;
        RECT 602.995 -23.965 603.325 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 -28.04 614.2 -27.72 ;
        RECT 612.515 -28.045 612.845 -27.715 ;
        RECT 611.155 -28.045 611.485 -27.715 ;
        RECT 609.795 -28.045 610.125 -27.715 ;
        RECT 608.435 -28.045 608.765 -27.715 ;
        RECT 604.355 -28.045 604.685 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 613.875 -34.845 614.205 -34.515 ;
        RECT 607.08 -34.84 614.205 -34.52 ;
        RECT 612.515 -34.845 612.845 -34.515 ;
        RECT 611.155 -34.845 611.485 -34.515 ;
        RECT 609.795 -34.845 610.125 -34.515 ;
        RECT 608.435 -34.845 608.765 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.08 -26.68 617.6 -26.36 ;
        RECT 615.235 -26.685 615.565 -26.355 ;
        RECT 612.515 -26.685 612.845 -26.355 ;
        RECT 611.155 -26.685 611.485 -26.355 ;
        RECT 609.795 -26.685 610.125 -26.355 ;
        RECT 608.435 -26.685 608.765 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.04 -29.4 628.48 -29.08 ;
        RECT 627.475 -29.405 627.805 -29.075 ;
        RECT 626.115 -29.405 626.445 -29.075 ;
        RECT 624.755 -29.405 625.085 -29.075 ;
        RECT 623.395 -29.405 623.725 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.28 -23.96 629.16 -23.64 ;
        RECT 627.475 -23.965 627.805 -23.635 ;
        RECT 626.115 -23.965 626.445 -23.635 ;
        RECT 624.755 -23.965 625.085 -23.635 ;
        RECT 623.395 -23.965 623.725 -23.635 ;
        RECT 622.035 -23.965 622.365 -23.635 ;
        RECT 619.315 -23.965 619.645 -23.635 ;
        RECT 617.955 -23.965 618.285 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.96 -28.04 629.16 -27.72 ;
        RECT 627.475 -28.045 627.805 -27.715 ;
        RECT 626.115 -28.045 626.445 -27.715 ;
        RECT 624.755 -28.045 625.085 -27.715 ;
        RECT 623.395 -28.045 623.725 -27.715 ;
        RECT 619.315 -28.045 619.645 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 628.835 -34.845 629.165 -34.515 ;
        RECT 622.04 -34.84 629.165 -34.52 ;
        RECT 627.475 -34.845 627.805 -34.515 ;
        RECT 626.115 -34.845 626.445 -34.515 ;
        RECT 624.755 -34.845 625.085 -34.515 ;
        RECT 623.395 -34.845 623.725 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.04 -26.68 632.56 -26.36 ;
        RECT 630.195 -26.685 630.525 -26.355 ;
        RECT 627.475 -26.685 627.805 -26.355 ;
        RECT 626.115 -26.685 626.445 -26.355 ;
        RECT 624.755 -26.685 625.085 -26.355 ;
        RECT 623.395 -26.685 623.725 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.24 -23.96 643.44 -23.64 ;
        RECT 641.075 -23.965 641.405 -23.635 ;
        RECT 639.715 -23.965 640.045 -23.635 ;
        RECT 638.355 -23.965 638.685 -23.635 ;
        RECT 636.995 -23.965 637.325 -23.635 ;
        RECT 634.275 -23.965 634.605 -23.635 ;
        RECT 632.915 -23.965 633.245 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.92 -28.04 643.44 -27.72 ;
        RECT 641.075 -28.045 641.405 -27.715 ;
        RECT 639.715 -28.045 640.045 -27.715 ;
        RECT 638.355 -28.045 638.685 -27.715 ;
        RECT 634.275 -28.045 634.605 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 637 -29.4 643.44 -29.08 ;
        RECT 641.075 -29.405 641.405 -29.075 ;
        RECT 639.715 -29.405 640.045 -29.075 ;
        RECT 638.355 -29.405 638.685 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 637 -34.84 643.44 -34.52 ;
        RECT 642.435 -34.845 642.765 -34.515 ;
        RECT 641.075 -34.845 641.405 -34.515 ;
        RECT 639.715 -34.845 640.045 -34.515 ;
        RECT 638.355 -34.845 638.685 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 637 -26.68 647.52 -26.36 ;
        RECT 645.155 -26.685 645.485 -26.355 ;
        RECT 641.075 -26.685 641.405 -26.355 ;
        RECT 639.715 -26.685 640.045 -26.355 ;
        RECT 638.355 -26.685 638.685 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.96 -29.4 657.72 -29.08 ;
        RECT 656.035 -29.405 656.365 -29.075 ;
        RECT 654.675 -29.405 655.005 -29.075 ;
        RECT 653.315 -29.405 653.645 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.2 -23.96 658.4 -23.64 ;
        RECT 656.035 -23.965 656.365 -23.635 ;
        RECT 654.675 -23.965 655.005 -23.635 ;
        RECT 653.315 -23.965 653.645 -23.635 ;
        RECT 651.955 -23.965 652.285 -23.635 ;
        RECT 649.235 -23.965 649.565 -23.635 ;
        RECT 647.875 -23.965 648.205 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.88 -28.04 658.4 -27.72 ;
        RECT 656.035 -28.045 656.365 -27.715 ;
        RECT 654.675 -28.045 655.005 -27.715 ;
        RECT 653.315 -28.045 653.645 -27.715 ;
        RECT 649.235 -28.045 649.565 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.96 -34.84 658.4 -34.52 ;
        RECT 657.395 -34.845 657.725 -34.515 ;
        RECT 656.035 -34.845 656.365 -34.515 ;
        RECT 654.675 -34.845 655.005 -34.515 ;
        RECT 653.315 -34.845 653.645 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.96 -26.68 662.48 -26.36 ;
        RECT 660.115 -26.685 660.445 -26.355 ;
        RECT 656.035 -26.685 656.365 -26.355 ;
        RECT 654.675 -26.685 655.005 -26.355 ;
        RECT 653.315 -26.685 653.645 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.92 -29.4 672.68 -29.08 ;
        RECT 670.995 -29.405 671.325 -29.075 ;
        RECT 669.635 -29.405 669.965 -29.075 ;
        RECT 668.275 -29.405 668.605 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.16 -23.96 673.36 -23.64 ;
        RECT 670.995 -23.965 671.325 -23.635 ;
        RECT 669.635 -23.965 669.965 -23.635 ;
        RECT 668.275 -23.965 668.605 -23.635 ;
        RECT 666.915 -23.965 667.245 -23.635 ;
        RECT 664.195 -23.965 664.525 -23.635 ;
        RECT 662.835 -23.965 663.165 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.84 -28.04 673.36 -27.72 ;
        RECT 670.995 -28.045 671.325 -27.715 ;
        RECT 669.635 -28.045 669.965 -27.715 ;
        RECT 668.275 -28.045 668.605 -27.715 ;
        RECT 664.195 -28.045 664.525 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.92 -34.84 673.36 -34.52 ;
        RECT 672.355 -34.845 672.685 -34.515 ;
        RECT 670.995 -34.845 671.325 -34.515 ;
        RECT 669.635 -34.845 669.965 -34.515 ;
        RECT 668.275 -34.845 668.605 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.92 -26.68 677.44 -26.36 ;
        RECT 675.075 -26.685 675.405 -26.355 ;
        RECT 670.995 -26.685 671.325 -26.355 ;
        RECT 669.635 -26.685 669.965 -26.355 ;
        RECT 668.275 -26.685 668.605 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 1.875 142.285 2.205 ;
        RECT 140.595 1.875 140.925 2.205 ;
        RECT 139.235 1.875 139.565 2.205 ;
        RECT 137.875 1.875 138.205 2.205 ;
        RECT 136.515 1.875 136.845 2.205 ;
        RECT 135.155 1.875 135.485 2.205 ;
        RECT 133.795 1.875 134.125 2.205 ;
        RECT 132.435 1.875 132.765 2.205 ;
        RECT 131.075 1.875 131.405 2.205 ;
        RECT 129.715 1.875 130.045 2.205 ;
        RECT 128.355 1.875 128.685 2.205 ;
        RECT 126.995 1.875 127.325 2.205 ;
        RECT 125.635 1.875 125.965 2.205 ;
        RECT 124.275 1.875 124.605 2.205 ;
        RECT 122.915 1.875 123.245 2.205 ;
        RECT 121.555 1.875 121.885 2.205 ;
        RECT 120.195 1.875 120.525 2.205 ;
        RECT 118.835 1.875 119.165 2.205 ;
        RECT 117.475 1.875 117.805 2.205 ;
        RECT 116.115 1.875 116.445 2.205 ;
        RECT 114.755 1.875 115.085 2.205 ;
        RECT 113.395 1.875 113.725 2.205 ;
        RECT 112.035 1.875 112.365 2.205 ;
        RECT 110.675 1.875 111.005 2.205 ;
        RECT 109.315 1.875 109.645 2.205 ;
        RECT 107.955 1.875 108.285 2.205 ;
        RECT 106.595 1.875 106.925 2.205 ;
        RECT 105.235 1.875 105.565 2.205 ;
        RECT 103.875 1.875 104.205 2.205 ;
        RECT 102.515 1.875 102.845 2.205 ;
        RECT 101.155 1.875 101.485 2.205 ;
        RECT 99.795 1.875 100.125 2.205 ;
        RECT 98.435 1.875 98.765 2.205 ;
        RECT 97.075 1.875 97.405 2.205 ;
        RECT 95.715 1.875 96.045 2.205 ;
        RECT 94.355 1.875 94.685 2.205 ;
        RECT 92.995 1.875 93.325 2.205 ;
        RECT 91.635 1.875 91.965 2.205 ;
        RECT 90.275 1.875 90.605 2.205 ;
        RECT 88.915 1.875 89.245 2.205 ;
        RECT 87.555 1.875 87.885 2.205 ;
        RECT 86.195 1.875 86.525 2.205 ;
        RECT 84.835 1.875 85.165 2.205 ;
        RECT 83.475 1.875 83.805 2.205 ;
        RECT 82.115 1.875 82.445 2.205 ;
        RECT 80.755 1.875 81.085 2.205 ;
        RECT 79.395 1.875 79.725 2.205 ;
        RECT 78.035 1.875 78.365 2.205 ;
        RECT 76.675 1.875 77.005 2.205 ;
        RECT 75.315 1.875 75.645 2.205 ;
        RECT 73.955 1.875 74.285 2.205 ;
        RECT 72.595 1.875 72.925 2.205 ;
        RECT 71.235 1.875 71.565 2.205 ;
        RECT 69.875 1.875 70.205 2.205 ;
        RECT 68.515 1.875 68.845 2.205 ;
        RECT 67.155 1.875 67.485 2.205 ;
        RECT 65.795 1.875 66.125 2.205 ;
        RECT 64.435 1.875 64.765 2.205 ;
        RECT 63.075 1.875 63.405 2.205 ;
        RECT 61.715 1.875 62.045 2.205 ;
        RECT 60.355 1.875 60.685 2.205 ;
        RECT 58.995 1.875 59.325 2.205 ;
        RECT 57.635 1.875 57.965 2.205 ;
        RECT 56.275 1.875 56.605 2.205 ;
        RECT 54.915 1.875 55.245 2.205 ;
        RECT 53.555 1.875 53.885 2.205 ;
        RECT 52.195 1.875 52.525 2.205 ;
        RECT 50.835 1.875 51.165 2.205 ;
        RECT 49.475 1.875 49.805 2.205 ;
        RECT 48.115 1.875 48.445 2.205 ;
        RECT 46.755 1.875 47.085 2.205 ;
        RECT 45.395 1.875 45.725 2.205 ;
        RECT 44.035 1.875 44.365 2.205 ;
        RECT 42.675 1.875 43.005 2.205 ;
        RECT 41.315 1.875 41.645 2.205 ;
        RECT 39.955 1.875 40.285 2.205 ;
        RECT 38.595 1.875 38.925 2.205 ;
        RECT 37.235 1.875 37.565 2.205 ;
        RECT 35.875 1.875 36.205 2.205 ;
        RECT 34.515 1.875 34.845 2.205 ;
        RECT 33.155 1.875 33.485 2.205 ;
        RECT 31.795 1.875 32.125 2.205 ;
        RECT 30.435 1.875 30.765 2.205 ;
        RECT 29.075 1.875 29.405 2.205 ;
        RECT 27.715 1.875 28.045 2.205 ;
        RECT 26.355 1.875 26.685 2.205 ;
        RECT 24.995 1.875 25.325 2.205 ;
        RECT 23.635 1.875 23.965 2.205 ;
        RECT 22.275 1.875 22.605 2.205 ;
        RECT 20.915 1.875 21.245 2.205 ;
        RECT 19.555 1.875 19.885 2.205 ;
        RECT 18.195 1.875 18.525 2.205 ;
        RECT 16.835 1.875 17.165 2.205 ;
        RECT 15.475 1.875 15.805 2.205 ;
        RECT 14.115 1.875 14.445 2.205 ;
        RECT 12.755 1.875 13.085 2.205 ;
        RECT 11.395 1.875 11.725 2.205 ;
        RECT 10.035 1.875 10.365 2.205 ;
        RECT 8.675 1.875 9.005 2.205 ;
        RECT 7.315 1.875 7.645 2.205 ;
        RECT 5.955 1.875 6.285 2.205 ;
        RECT 4.595 1.875 4.925 2.205 ;
        RECT 3.235 1.875 3.565 2.205 ;
        RECT 1.875 1.875 2.205 2.205 ;
        RECT 0.515 1.875 0.845 2.205 ;
        RECT -0.845 1.875 -0.515 2.205 ;
        RECT 677.795 1.875 678.125 2.205 ;
        RECT -1.52 1.88 678.125 2.2 ;
        RECT 676.435 1.875 676.765 2.205 ;
        RECT 675.075 1.875 675.405 2.205 ;
        RECT 673.715 1.875 674.045 2.205 ;
        RECT 672.355 1.875 672.685 2.205 ;
        RECT 670.995 1.875 671.325 2.205 ;
        RECT 669.635 1.875 669.965 2.205 ;
        RECT 668.275 1.875 668.605 2.205 ;
        RECT 666.915 1.875 667.245 2.205 ;
        RECT 665.555 1.875 665.885 2.205 ;
        RECT 664.195 1.875 664.525 2.205 ;
        RECT 662.835 1.875 663.165 2.205 ;
        RECT 661.475 1.875 661.805 2.205 ;
        RECT 660.115 1.875 660.445 2.205 ;
        RECT 658.755 1.875 659.085 2.205 ;
        RECT 657.395 1.875 657.725 2.205 ;
        RECT 656.035 1.875 656.365 2.205 ;
        RECT 654.675 1.875 655.005 2.205 ;
        RECT 653.315 1.875 653.645 2.205 ;
        RECT 651.955 1.875 652.285 2.205 ;
        RECT 650.595 1.875 650.925 2.205 ;
        RECT 649.235 1.875 649.565 2.205 ;
        RECT 647.875 1.875 648.205 2.205 ;
        RECT 646.515 1.875 646.845 2.205 ;
        RECT 645.155 1.875 645.485 2.205 ;
        RECT 643.795 1.875 644.125 2.205 ;
        RECT 642.435 1.875 642.765 2.205 ;
        RECT 641.075 1.875 641.405 2.205 ;
        RECT 639.715 1.875 640.045 2.205 ;
        RECT 638.355 1.875 638.685 2.205 ;
        RECT 636.995 1.875 637.325 2.205 ;
        RECT 635.635 1.875 635.965 2.205 ;
        RECT 634.275 1.875 634.605 2.205 ;
        RECT 632.915 1.875 633.245 2.205 ;
        RECT 631.555 1.875 631.885 2.205 ;
        RECT 630.195 1.875 630.525 2.205 ;
        RECT 628.835 1.875 629.165 2.205 ;
        RECT 627.475 1.875 627.805 2.205 ;
        RECT 626.115 1.875 626.445 2.205 ;
        RECT 624.755 1.875 625.085 2.205 ;
        RECT 623.395 1.875 623.725 2.205 ;
        RECT 622.035 1.875 622.365 2.205 ;
        RECT 620.675 1.875 621.005 2.205 ;
        RECT 619.315 1.875 619.645 2.205 ;
        RECT 617.955 1.875 618.285 2.205 ;
        RECT 616.595 1.875 616.925 2.205 ;
        RECT 615.235 1.875 615.565 2.205 ;
        RECT 613.875 1.875 614.205 2.205 ;
        RECT 612.515 1.875 612.845 2.205 ;
        RECT 611.155 1.875 611.485 2.205 ;
        RECT 609.795 1.875 610.125 2.205 ;
        RECT 608.435 1.875 608.765 2.205 ;
        RECT 607.075 1.875 607.405 2.205 ;
        RECT 605.715 1.875 606.045 2.205 ;
        RECT 604.355 1.875 604.685 2.205 ;
        RECT 602.995 1.875 603.325 2.205 ;
        RECT 601.635 1.875 601.965 2.205 ;
        RECT 600.275 1.875 600.605 2.205 ;
        RECT 598.915 1.875 599.245 2.205 ;
        RECT 597.555 1.875 597.885 2.205 ;
        RECT 596.195 1.875 596.525 2.205 ;
        RECT 594.835 1.875 595.165 2.205 ;
        RECT 593.475 1.875 593.805 2.205 ;
        RECT 592.115 1.875 592.445 2.205 ;
        RECT 590.755 1.875 591.085 2.205 ;
        RECT 589.395 1.875 589.725 2.205 ;
        RECT 588.035 1.875 588.365 2.205 ;
        RECT 586.675 1.875 587.005 2.205 ;
        RECT 585.315 1.875 585.645 2.205 ;
        RECT 583.955 1.875 584.285 2.205 ;
        RECT 582.595 1.875 582.925 2.205 ;
        RECT 581.235 1.875 581.565 2.205 ;
        RECT 579.875 1.875 580.205 2.205 ;
        RECT 578.515 1.875 578.845 2.205 ;
        RECT 577.155 1.875 577.485 2.205 ;
        RECT 575.795 1.875 576.125 2.205 ;
        RECT 574.435 1.875 574.765 2.205 ;
        RECT 573.075 1.875 573.405 2.205 ;
        RECT 571.715 1.875 572.045 2.205 ;
        RECT 570.355 1.875 570.685 2.205 ;
        RECT 568.995 1.875 569.325 2.205 ;
        RECT 567.635 1.875 567.965 2.205 ;
        RECT 566.275 1.875 566.605 2.205 ;
        RECT 564.915 1.875 565.245 2.205 ;
        RECT 563.555 1.875 563.885 2.205 ;
        RECT 562.195 1.875 562.525 2.205 ;
        RECT 560.835 1.875 561.165 2.205 ;
        RECT 559.475 1.875 559.805 2.205 ;
        RECT 558.115 1.875 558.445 2.205 ;
        RECT 556.755 1.875 557.085 2.205 ;
        RECT 555.395 1.875 555.725 2.205 ;
        RECT 554.035 1.875 554.365 2.205 ;
        RECT 552.675 1.875 553.005 2.205 ;
        RECT 551.315 1.875 551.645 2.205 ;
        RECT 549.955 1.875 550.285 2.205 ;
        RECT 548.595 1.875 548.925 2.205 ;
        RECT 547.235 1.875 547.565 2.205 ;
        RECT 545.875 1.875 546.205 2.205 ;
        RECT 544.515 1.875 544.845 2.205 ;
        RECT 543.155 1.875 543.485 2.205 ;
        RECT 541.795 1.875 542.125 2.205 ;
        RECT 540.435 1.875 540.765 2.205 ;
        RECT 539.075 1.875 539.405 2.205 ;
        RECT 537.715 1.875 538.045 2.205 ;
        RECT 536.355 1.875 536.685 2.205 ;
        RECT 534.995 1.875 535.325 2.205 ;
        RECT 533.635 1.875 533.965 2.205 ;
        RECT 532.275 1.875 532.605 2.205 ;
        RECT 530.915 1.875 531.245 2.205 ;
        RECT 529.555 1.875 529.885 2.205 ;
        RECT 528.195 1.875 528.525 2.205 ;
        RECT 526.835 1.875 527.165 2.205 ;
        RECT 525.475 1.875 525.805 2.205 ;
        RECT 524.115 1.875 524.445 2.205 ;
        RECT 522.755 1.875 523.085 2.205 ;
        RECT 521.395 1.875 521.725 2.205 ;
        RECT 520.035 1.875 520.365 2.205 ;
        RECT 518.675 1.875 519.005 2.205 ;
        RECT 517.315 1.875 517.645 2.205 ;
        RECT 515.955 1.875 516.285 2.205 ;
        RECT 514.595 1.875 514.925 2.205 ;
        RECT 513.235 1.875 513.565 2.205 ;
        RECT 511.875 1.875 512.205 2.205 ;
        RECT 510.515 1.875 510.845 2.205 ;
        RECT 509.155 1.875 509.485 2.205 ;
        RECT 507.795 1.875 508.125 2.205 ;
        RECT 506.435 1.875 506.765 2.205 ;
        RECT 505.075 1.875 505.405 2.205 ;
        RECT 503.715 1.875 504.045 2.205 ;
        RECT 502.355 1.875 502.685 2.205 ;
        RECT 500.995 1.875 501.325 2.205 ;
        RECT 499.635 1.875 499.965 2.205 ;
        RECT 498.275 1.875 498.605 2.205 ;
        RECT 496.915 1.875 497.245 2.205 ;
        RECT 495.555 1.875 495.885 2.205 ;
        RECT 494.195 1.875 494.525 2.205 ;
        RECT 492.835 1.875 493.165 2.205 ;
        RECT 491.475 1.875 491.805 2.205 ;
        RECT 490.115 1.875 490.445 2.205 ;
        RECT 488.755 1.875 489.085 2.205 ;
        RECT 487.395 1.875 487.725 2.205 ;
        RECT 486.035 1.875 486.365 2.205 ;
        RECT 484.675 1.875 485.005 2.205 ;
        RECT 483.315 1.875 483.645 2.205 ;
        RECT 481.955 1.875 482.285 2.205 ;
        RECT 480.595 1.875 480.925 2.205 ;
        RECT 479.235 1.875 479.565 2.205 ;
        RECT 477.875 1.875 478.205 2.205 ;
        RECT 476.515 1.875 476.845 2.205 ;
        RECT 475.155 1.875 475.485 2.205 ;
        RECT 473.795 1.875 474.125 2.205 ;
        RECT 472.435 1.875 472.765 2.205 ;
        RECT 471.075 1.875 471.405 2.205 ;
        RECT 469.715 1.875 470.045 2.205 ;
        RECT 468.355 1.875 468.685 2.205 ;
        RECT 466.995 1.875 467.325 2.205 ;
        RECT 465.635 1.875 465.965 2.205 ;
        RECT 464.275 1.875 464.605 2.205 ;
        RECT 462.915 1.875 463.245 2.205 ;
        RECT 461.555 1.875 461.885 2.205 ;
        RECT 460.195 1.875 460.525 2.205 ;
        RECT 458.835 1.875 459.165 2.205 ;
        RECT 457.475 1.875 457.805 2.205 ;
        RECT 456.115 1.875 456.445 2.205 ;
        RECT 454.755 1.875 455.085 2.205 ;
        RECT 453.395 1.875 453.725 2.205 ;
        RECT 452.035 1.875 452.365 2.205 ;
        RECT 450.675 1.875 451.005 2.205 ;
        RECT 449.315 1.875 449.645 2.205 ;
        RECT 447.955 1.875 448.285 2.205 ;
        RECT 446.595 1.875 446.925 2.205 ;
        RECT 445.235 1.875 445.565 2.205 ;
        RECT 443.875 1.875 444.205 2.205 ;
        RECT 442.515 1.875 442.845 2.205 ;
        RECT 441.155 1.875 441.485 2.205 ;
        RECT 439.795 1.875 440.125 2.205 ;
        RECT 438.435 1.875 438.765 2.205 ;
        RECT 437.075 1.875 437.405 2.205 ;
        RECT 435.715 1.875 436.045 2.205 ;
        RECT 434.355 1.875 434.685 2.205 ;
        RECT 432.995 1.875 433.325 2.205 ;
        RECT 431.635 1.875 431.965 2.205 ;
        RECT 430.275 1.875 430.605 2.205 ;
        RECT 428.915 1.875 429.245 2.205 ;
        RECT 427.555 1.875 427.885 2.205 ;
        RECT 426.195 1.875 426.525 2.205 ;
        RECT 424.835 1.875 425.165 2.205 ;
        RECT 423.475 1.875 423.805 2.205 ;
        RECT 422.115 1.875 422.445 2.205 ;
        RECT 420.755 1.875 421.085 2.205 ;
        RECT 419.395 1.875 419.725 2.205 ;
        RECT 418.035 1.875 418.365 2.205 ;
        RECT 416.675 1.875 417.005 2.205 ;
        RECT 415.315 1.875 415.645 2.205 ;
        RECT 413.955 1.875 414.285 2.205 ;
        RECT 412.595 1.875 412.925 2.205 ;
        RECT 411.235 1.875 411.565 2.205 ;
        RECT 409.875 1.875 410.205 2.205 ;
        RECT 408.515 1.875 408.845 2.205 ;
        RECT 407.155 1.875 407.485 2.205 ;
        RECT 405.795 1.875 406.125 2.205 ;
        RECT 404.435 1.875 404.765 2.205 ;
        RECT 403.075 1.875 403.405 2.205 ;
        RECT 401.715 1.875 402.045 2.205 ;
        RECT 400.355 1.875 400.685 2.205 ;
        RECT 398.995 1.875 399.325 2.205 ;
        RECT 397.635 1.875 397.965 2.205 ;
        RECT 396.275 1.875 396.605 2.205 ;
        RECT 394.915 1.875 395.245 2.205 ;
        RECT 393.555 1.875 393.885 2.205 ;
        RECT 392.195 1.875 392.525 2.205 ;
        RECT 390.835 1.875 391.165 2.205 ;
        RECT 389.475 1.875 389.805 2.205 ;
        RECT 388.115 1.875 388.445 2.205 ;
        RECT 386.755 1.875 387.085 2.205 ;
        RECT 385.395 1.875 385.725 2.205 ;
        RECT 384.035 1.875 384.365 2.205 ;
        RECT 382.675 1.875 383.005 2.205 ;
        RECT 381.315 1.875 381.645 2.205 ;
        RECT 379.955 1.875 380.285 2.205 ;
        RECT 378.595 1.875 378.925 2.205 ;
        RECT 377.235 1.875 377.565 2.205 ;
        RECT 375.875 1.875 376.205 2.205 ;
        RECT 374.515 1.875 374.845 2.205 ;
        RECT 373.155 1.875 373.485 2.205 ;
        RECT 371.795 1.875 372.125 2.205 ;
        RECT 370.435 1.875 370.765 2.205 ;
        RECT 369.075 1.875 369.405 2.205 ;
        RECT 367.715 1.875 368.045 2.205 ;
        RECT 366.355 1.875 366.685 2.205 ;
        RECT 364.995 1.875 365.325 2.205 ;
        RECT 363.635 1.875 363.965 2.205 ;
        RECT 362.275 1.875 362.605 2.205 ;
        RECT 360.915 1.875 361.245 2.205 ;
        RECT 359.555 1.875 359.885 2.205 ;
        RECT 358.195 1.875 358.525 2.205 ;
        RECT 356.835 1.875 357.165 2.205 ;
        RECT 355.475 1.875 355.805 2.205 ;
        RECT 354.115 1.875 354.445 2.205 ;
        RECT 352.755 1.875 353.085 2.205 ;
        RECT 351.395 1.875 351.725 2.205 ;
        RECT 350.035 1.875 350.365 2.205 ;
        RECT 348.675 1.875 349.005 2.205 ;
        RECT 347.315 1.875 347.645 2.205 ;
        RECT 345.955 1.875 346.285 2.205 ;
        RECT 344.595 1.875 344.925 2.205 ;
        RECT 343.235 1.875 343.565 2.205 ;
        RECT 341.875 1.875 342.205 2.205 ;
        RECT 340.515 1.875 340.845 2.205 ;
        RECT 339.155 1.875 339.485 2.205 ;
        RECT 337.795 1.875 338.125 2.205 ;
        RECT 336.435 1.875 336.765 2.205 ;
        RECT 335.075 1.875 335.405 2.205 ;
        RECT 333.715 1.875 334.045 2.205 ;
        RECT 332.355 1.875 332.685 2.205 ;
        RECT 330.995 1.875 331.325 2.205 ;
        RECT 329.635 1.875 329.965 2.205 ;
        RECT 328.275 1.875 328.605 2.205 ;
        RECT 326.915 1.875 327.245 2.205 ;
        RECT 325.555 1.875 325.885 2.205 ;
        RECT 324.195 1.875 324.525 2.205 ;
        RECT 322.835 1.875 323.165 2.205 ;
        RECT 321.475 1.875 321.805 2.205 ;
        RECT 320.115 1.875 320.445 2.205 ;
        RECT 318.755 1.875 319.085 2.205 ;
        RECT 317.395 1.875 317.725 2.205 ;
        RECT 316.035 1.875 316.365 2.205 ;
        RECT 314.675 1.875 315.005 2.205 ;
        RECT 313.315 1.875 313.645 2.205 ;
        RECT 311.955 1.875 312.285 2.205 ;
        RECT 310.595 1.875 310.925 2.205 ;
        RECT 309.235 1.875 309.565 2.205 ;
        RECT 307.875 1.875 308.205 2.205 ;
        RECT 306.515 1.875 306.845 2.205 ;
        RECT 305.155 1.875 305.485 2.205 ;
        RECT 303.795 1.875 304.125 2.205 ;
        RECT 302.435 1.875 302.765 2.205 ;
        RECT 301.075 1.875 301.405 2.205 ;
        RECT 299.715 1.875 300.045 2.205 ;
        RECT 298.355 1.875 298.685 2.205 ;
        RECT 296.995 1.875 297.325 2.205 ;
        RECT 295.635 1.875 295.965 2.205 ;
        RECT 294.275 1.875 294.605 2.205 ;
        RECT 292.915 1.875 293.245 2.205 ;
        RECT 291.555 1.875 291.885 2.205 ;
        RECT 290.195 1.875 290.525 2.205 ;
        RECT 288.835 1.875 289.165 2.205 ;
        RECT 287.475 1.875 287.805 2.205 ;
        RECT 286.115 1.875 286.445 2.205 ;
        RECT 284.755 1.875 285.085 2.205 ;
        RECT 283.395 1.875 283.725 2.205 ;
        RECT 282.035 1.875 282.365 2.205 ;
        RECT 280.675 1.875 281.005 2.205 ;
        RECT 279.315 1.875 279.645 2.205 ;
        RECT 277.955 1.875 278.285 2.205 ;
        RECT 276.595 1.875 276.925 2.205 ;
        RECT 275.235 1.875 275.565 2.205 ;
        RECT 273.875 1.875 274.205 2.205 ;
        RECT 272.515 1.875 272.845 2.205 ;
        RECT 271.155 1.875 271.485 2.205 ;
        RECT 269.795 1.875 270.125 2.205 ;
        RECT 268.435 1.875 268.765 2.205 ;
        RECT 267.075 1.875 267.405 2.205 ;
        RECT 265.715 1.875 266.045 2.205 ;
        RECT 264.355 1.875 264.685 2.205 ;
        RECT 262.995 1.875 263.325 2.205 ;
        RECT 261.635 1.875 261.965 2.205 ;
        RECT 260.275 1.875 260.605 2.205 ;
        RECT 258.915 1.875 259.245 2.205 ;
        RECT 257.555 1.875 257.885 2.205 ;
        RECT 256.195 1.875 256.525 2.205 ;
        RECT 254.835 1.875 255.165 2.205 ;
        RECT 253.475 1.875 253.805 2.205 ;
        RECT 252.115 1.875 252.445 2.205 ;
        RECT 250.755 1.875 251.085 2.205 ;
        RECT 249.395 1.875 249.725 2.205 ;
        RECT 248.035 1.875 248.365 2.205 ;
        RECT 246.675 1.875 247.005 2.205 ;
        RECT 245.315 1.875 245.645 2.205 ;
        RECT 243.955 1.875 244.285 2.205 ;
        RECT 242.595 1.875 242.925 2.205 ;
        RECT 241.235 1.875 241.565 2.205 ;
        RECT 239.875 1.875 240.205 2.205 ;
        RECT 238.515 1.875 238.845 2.205 ;
        RECT 237.155 1.875 237.485 2.205 ;
        RECT 235.795 1.875 236.125 2.205 ;
        RECT 234.435 1.875 234.765 2.205 ;
        RECT 233.075 1.875 233.405 2.205 ;
        RECT 231.715 1.875 232.045 2.205 ;
        RECT 230.355 1.875 230.685 2.205 ;
        RECT 228.995 1.875 229.325 2.205 ;
        RECT 227.635 1.875 227.965 2.205 ;
        RECT 226.275 1.875 226.605 2.205 ;
        RECT 224.915 1.875 225.245 2.205 ;
        RECT 223.555 1.875 223.885 2.205 ;
        RECT 222.195 1.875 222.525 2.205 ;
        RECT 220.835 1.875 221.165 2.205 ;
        RECT 219.475 1.875 219.805 2.205 ;
        RECT 218.115 1.875 218.445 2.205 ;
        RECT 216.755 1.875 217.085 2.205 ;
        RECT 215.395 1.875 215.725 2.205 ;
        RECT 214.035 1.875 214.365 2.205 ;
        RECT 212.675 1.875 213.005 2.205 ;
        RECT 211.315 1.875 211.645 2.205 ;
        RECT 209.955 1.875 210.285 2.205 ;
        RECT 208.595 1.875 208.925 2.205 ;
        RECT 207.235 1.875 207.565 2.205 ;
        RECT 205.875 1.875 206.205 2.205 ;
        RECT 204.515 1.875 204.845 2.205 ;
        RECT 203.155 1.875 203.485 2.205 ;
        RECT 201.795 1.875 202.125 2.205 ;
        RECT 200.435 1.875 200.765 2.205 ;
        RECT 199.075 1.875 199.405 2.205 ;
        RECT 197.715 1.875 198.045 2.205 ;
        RECT 196.355 1.875 196.685 2.205 ;
        RECT 194.995 1.875 195.325 2.205 ;
        RECT 193.635 1.875 193.965 2.205 ;
        RECT 192.275 1.875 192.605 2.205 ;
        RECT 190.915 1.875 191.245 2.205 ;
        RECT 189.555 1.875 189.885 2.205 ;
        RECT 188.195 1.875 188.525 2.205 ;
        RECT 186.835 1.875 187.165 2.205 ;
        RECT 185.475 1.875 185.805 2.205 ;
        RECT 184.115 1.875 184.445 2.205 ;
        RECT 182.755 1.875 183.085 2.205 ;
        RECT 181.395 1.875 181.725 2.205 ;
        RECT 180.035 1.875 180.365 2.205 ;
        RECT 178.675 1.875 179.005 2.205 ;
        RECT 177.315 1.875 177.645 2.205 ;
        RECT 175.955 1.875 176.285 2.205 ;
        RECT 174.595 1.875 174.925 2.205 ;
        RECT 173.235 1.875 173.565 2.205 ;
        RECT 171.875 1.875 172.205 2.205 ;
        RECT 170.515 1.875 170.845 2.205 ;
        RECT 169.155 1.875 169.485 2.205 ;
        RECT 167.795 1.875 168.125 2.205 ;
        RECT 166.435 1.875 166.765 2.205 ;
        RECT 165.075 1.875 165.405 2.205 ;
        RECT 163.715 1.875 164.045 2.205 ;
        RECT 162.355 1.875 162.685 2.205 ;
        RECT 160.995 1.875 161.325 2.205 ;
        RECT 159.635 1.875 159.965 2.205 ;
        RECT 158.275 1.875 158.605 2.205 ;
        RECT 156.915 1.875 157.245 2.205 ;
        RECT 155.555 1.875 155.885 2.205 ;
        RECT 154.195 1.875 154.525 2.205 ;
        RECT 152.835 1.875 153.165 2.205 ;
        RECT 151.475 1.875 151.805 2.205 ;
        RECT 150.115 1.875 150.445 2.205 ;
        RECT 148.755 1.875 149.085 2.205 ;
        RECT 147.395 1.875 147.725 2.205 ;
        RECT 146.035 1.875 146.365 2.205 ;
        RECT 144.675 1.875 145.005 2.205 ;
        RECT 143.315 1.875 143.645 2.205 ;
        RECT 789.315 1.875 789.645 2.205 ;
        RECT 787.955 1.875 788.285 2.205 ;
        RECT 786.595 1.875 786.925 2.205 ;
        RECT 785.235 1.875 785.565 2.205 ;
        RECT 783.875 1.875 784.205 2.205 ;
        RECT 782.515 1.875 782.845 2.205 ;
        RECT 781.155 1.875 781.485 2.205 ;
        RECT 779.795 1.875 780.125 2.205 ;
        RECT 778.435 1.875 778.765 2.205 ;
        RECT 777.075 1.875 777.405 2.205 ;
        RECT 775.715 1.875 776.045 2.205 ;
        RECT 774.355 1.875 774.685 2.205 ;
        RECT 772.995 1.875 773.325 2.205 ;
        RECT 771.635 1.875 771.965 2.205 ;
        RECT 770.275 1.875 770.605 2.205 ;
        RECT 768.915 1.875 769.245 2.205 ;
        RECT 767.555 1.875 767.885 2.205 ;
        RECT 766.195 1.875 766.525 2.205 ;
        RECT 764.835 1.875 765.165 2.205 ;
        RECT 763.475 1.875 763.805 2.205 ;
        RECT 762.115 1.875 762.445 2.205 ;
        RECT 760.755 1.875 761.085 2.205 ;
        RECT 759.395 1.875 759.725 2.205 ;
        RECT 758.035 1.875 758.365 2.205 ;
        RECT 756.675 1.875 757.005 2.205 ;
        RECT 755.315 1.875 755.645 2.205 ;
        RECT 753.955 1.875 754.285 2.205 ;
        RECT 752.595 1.875 752.925 2.205 ;
        RECT 751.235 1.875 751.565 2.205 ;
        RECT 749.875 1.875 750.205 2.205 ;
        RECT 748.515 1.875 748.845 2.205 ;
        RECT 747.155 1.875 747.485 2.205 ;
        RECT 745.795 1.875 746.125 2.205 ;
        RECT 744.435 1.875 744.765 2.205 ;
        RECT 743.075 1.875 743.405 2.205 ;
        RECT 741.715 1.875 742.045 2.205 ;
        RECT 740.355 1.875 740.685 2.205 ;
        RECT 738.995 1.875 739.325 2.205 ;
        RECT 737.635 1.875 737.965 2.205 ;
        RECT 736.275 1.875 736.605 2.205 ;
        RECT 734.915 1.875 735.245 2.205 ;
        RECT 733.555 1.875 733.885 2.205 ;
        RECT 732.195 1.875 732.525 2.205 ;
        RECT 730.835 1.875 731.165 2.205 ;
        RECT 729.475 1.875 729.805 2.205 ;
        RECT 728.115 1.875 728.445 2.205 ;
        RECT 726.755 1.875 727.085 2.205 ;
        RECT 725.395 1.875 725.725 2.205 ;
        RECT 724.035 1.875 724.365 2.205 ;
        RECT 722.675 1.875 723.005 2.205 ;
        RECT 721.315 1.875 721.645 2.205 ;
        RECT 719.955 1.875 720.285 2.205 ;
        RECT 718.595 1.875 718.925 2.205 ;
        RECT 717.235 1.875 717.565 2.205 ;
        RECT 715.875 1.875 716.205 2.205 ;
        RECT 714.515 1.875 714.845 2.205 ;
        RECT 713.155 1.875 713.485 2.205 ;
        RECT 711.795 1.875 712.125 2.205 ;
        RECT 710.435 1.875 710.765 2.205 ;
        RECT 709.075 1.875 709.405 2.205 ;
        RECT 707.715 1.875 708.045 2.205 ;
        RECT 706.355 1.875 706.685 2.205 ;
        RECT 704.995 1.875 705.325 2.205 ;
        RECT 703.635 1.875 703.965 2.205 ;
        RECT 702.275 1.875 702.605 2.205 ;
        RECT 700.915 1.875 701.245 2.205 ;
        RECT 699.555 1.875 699.885 2.205 ;
        RECT 698.195 1.875 698.525 2.205 ;
        RECT 696.835 1.875 697.165 2.205 ;
        RECT 695.475 1.875 695.805 2.205 ;
        RECT 694.115 1.875 694.445 2.205 ;
        RECT 692.755 1.875 693.085 2.205 ;
        RECT 691.395 1.875 691.725 2.205 ;
        RECT 690.035 1.875 690.365 2.205 ;
        RECT 688.675 1.875 689.005 2.205 ;
        RECT 687.315 1.875 687.645 2.205 ;
        RECT 685.955 1.875 686.285 2.205 ;
        RECT 684.595 1.875 684.925 2.205 ;
        RECT 683.235 1.875 683.565 2.205 ;
        RECT 681.875 1.875 682.205 2.205 ;
        RECT 680.515 1.875 680.845 2.205 ;
        RECT 679.155 1.875 679.485 2.205 ;
        RECT 678.125 1.88 954.88 2.2 ;
        RECT 953.875 1.875 954.205 2.205 ;
        RECT 952.515 1.875 952.845 2.205 ;
        RECT 951.155 1.875 951.485 2.205 ;
        RECT 949.795 1.875 950.125 2.205 ;
        RECT 948.435 1.875 948.765 2.205 ;
        RECT 947.075 1.875 947.405 2.205 ;
        RECT 945.715 1.875 946.045 2.205 ;
        RECT 944.355 1.875 944.685 2.205 ;
        RECT 942.995 1.875 943.325 2.205 ;
        RECT 941.635 1.875 941.965 2.205 ;
        RECT 940.275 1.875 940.605 2.205 ;
        RECT 938.915 1.875 939.245 2.205 ;
        RECT 937.555 1.875 937.885 2.205 ;
        RECT 936.195 1.875 936.525 2.205 ;
        RECT 934.835 1.875 935.165 2.205 ;
        RECT 933.475 1.875 933.805 2.205 ;
        RECT 932.115 1.875 932.445 2.205 ;
        RECT 930.755 1.875 931.085 2.205 ;
        RECT 929.395 1.875 929.725 2.205 ;
        RECT 928.035 1.875 928.365 2.205 ;
        RECT 926.675 1.875 927.005 2.205 ;
        RECT 925.315 1.875 925.645 2.205 ;
        RECT 923.955 1.875 924.285 2.205 ;
        RECT 922.595 1.875 922.925 2.205 ;
        RECT 921.235 1.875 921.565 2.205 ;
        RECT 919.875 1.875 920.205 2.205 ;
        RECT 918.515 1.875 918.845 2.205 ;
        RECT 917.155 1.875 917.485 2.205 ;
        RECT 915.795 1.875 916.125 2.205 ;
        RECT 914.435 1.875 914.765 2.205 ;
        RECT 913.075 1.875 913.405 2.205 ;
        RECT 911.715 1.875 912.045 2.205 ;
        RECT 910.355 1.875 910.685 2.205 ;
        RECT 908.995 1.875 909.325 2.205 ;
        RECT 907.635 1.875 907.965 2.205 ;
        RECT 906.275 1.875 906.605 2.205 ;
        RECT 904.915 1.875 905.245 2.205 ;
        RECT 903.555 1.875 903.885 2.205 ;
        RECT 902.195 1.875 902.525 2.205 ;
        RECT 900.835 1.875 901.165 2.205 ;
        RECT 899.475 1.875 899.805 2.205 ;
        RECT 898.115 1.875 898.445 2.205 ;
        RECT 896.755 1.875 897.085 2.205 ;
        RECT 895.395 1.875 895.725 2.205 ;
        RECT 894.035 1.875 894.365 2.205 ;
        RECT 892.675 1.875 893.005 2.205 ;
        RECT 891.315 1.875 891.645 2.205 ;
        RECT 889.955 1.875 890.285 2.205 ;
        RECT 888.595 1.875 888.925 2.205 ;
        RECT 887.235 1.875 887.565 2.205 ;
        RECT 885.875 1.875 886.205 2.205 ;
        RECT 884.515 1.875 884.845 2.205 ;
        RECT 883.155 1.875 883.485 2.205 ;
        RECT 881.795 1.875 882.125 2.205 ;
        RECT 880.435 1.875 880.765 2.205 ;
        RECT 879.075 1.875 879.405 2.205 ;
        RECT 877.715 1.875 878.045 2.205 ;
        RECT 876.355 1.875 876.685 2.205 ;
        RECT 874.995 1.875 875.325 2.205 ;
        RECT 873.635 1.875 873.965 2.205 ;
        RECT 872.275 1.875 872.605 2.205 ;
        RECT 870.915 1.875 871.245 2.205 ;
        RECT 869.555 1.875 869.885 2.205 ;
        RECT 868.195 1.875 868.525 2.205 ;
        RECT 866.835 1.875 867.165 2.205 ;
        RECT 865.475 1.875 865.805 2.205 ;
        RECT 864.115 1.875 864.445 2.205 ;
        RECT 862.755 1.875 863.085 2.205 ;
        RECT 861.395 1.875 861.725 2.205 ;
        RECT 860.035 1.875 860.365 2.205 ;
        RECT 858.675 1.875 859.005 2.205 ;
        RECT 857.315 1.875 857.645 2.205 ;
        RECT 855.955 1.875 856.285 2.205 ;
        RECT 854.595 1.875 854.925 2.205 ;
        RECT 853.235 1.875 853.565 2.205 ;
        RECT 851.875 1.875 852.205 2.205 ;
        RECT 850.515 1.875 850.845 2.205 ;
        RECT 849.155 1.875 849.485 2.205 ;
        RECT 847.795 1.875 848.125 2.205 ;
        RECT 846.435 1.875 846.765 2.205 ;
        RECT 845.075 1.875 845.405 2.205 ;
        RECT 843.715 1.875 844.045 2.205 ;
        RECT 842.355 1.875 842.685 2.205 ;
        RECT 840.995 1.875 841.325 2.205 ;
        RECT 839.635 1.875 839.965 2.205 ;
        RECT 838.275 1.875 838.605 2.205 ;
        RECT 836.915 1.875 837.245 2.205 ;
        RECT 835.555 1.875 835.885 2.205 ;
        RECT 834.195 1.875 834.525 2.205 ;
        RECT 832.835 1.875 833.165 2.205 ;
        RECT 831.475 1.875 831.805 2.205 ;
        RECT 830.115 1.875 830.445 2.205 ;
        RECT 828.755 1.875 829.085 2.205 ;
        RECT 827.395 1.875 827.725 2.205 ;
        RECT 826.035 1.875 826.365 2.205 ;
        RECT 824.675 1.875 825.005 2.205 ;
        RECT 823.315 1.875 823.645 2.205 ;
        RECT 821.955 1.875 822.285 2.205 ;
        RECT 820.595 1.875 820.925 2.205 ;
        RECT 819.235 1.875 819.565 2.205 ;
        RECT 817.875 1.875 818.205 2.205 ;
        RECT 816.515 1.875 816.845 2.205 ;
        RECT 815.155 1.875 815.485 2.205 ;
        RECT 813.795 1.875 814.125 2.205 ;
        RECT 812.435 1.875 812.765 2.205 ;
        RECT 811.075 1.875 811.405 2.205 ;
        RECT 809.715 1.875 810.045 2.205 ;
        RECT 808.355 1.875 808.685 2.205 ;
        RECT 806.995 1.875 807.325 2.205 ;
        RECT 805.635 1.875 805.965 2.205 ;
        RECT 804.275 1.875 804.605 2.205 ;
        RECT 802.915 1.875 803.245 2.205 ;
        RECT 801.555 1.875 801.885 2.205 ;
        RECT 800.195 1.875 800.525 2.205 ;
        RECT 798.835 1.875 799.165 2.205 ;
        RECT 797.475 1.875 797.805 2.205 ;
        RECT 796.115 1.875 796.445 2.205 ;
        RECT 794.755 1.875 795.085 2.205 ;
        RECT 793.395 1.875 793.725 2.205 ;
        RECT 792.035 1.875 792.365 2.205 ;
        RECT 790.675 1.875 791.005 2.205 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -23.96 2.88 -23.64 ;
        RECT 0.515 -23.965 0.845 -23.635 ;
        RECT -0.845 -23.965 -0.515 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -34.84 5.6 -34.52 ;
        RECT 4.595 -34.845 4.925 -34.515 ;
        RECT 3.235 -34.845 3.565 -34.515 ;
        RECT 1.875 -34.845 2.205 -34.515 ;
        RECT 0.515 -34.845 0.845 -34.515 ;
        RECT -0.845 -34.845 -0.515 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -29.4 17.16 -29.08 ;
        RECT 15.475 -29.405 15.805 -29.075 ;
        RECT 14.115 -29.405 14.445 -29.075 ;
        RECT 12.755 -29.405 13.085 -29.075 ;
        RECT 11.395 -29.405 11.725 -29.075 ;
        RECT 8.675 -29.405 9.005 -29.075 ;
        RECT 7.315 -29.405 7.645 -29.075 ;
        RECT 5.955 -29.405 6.285 -29.075 ;
        RECT 4.595 -29.405 4.925 -29.075 ;
        RECT 3.235 -29.405 3.565 -29.075 ;
        RECT 1.875 -29.405 2.205 -29.075 ;
        RECT 0.515 -29.405 0.845 -29.075 ;
        RECT -0.845 -29.405 -0.515 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.64 -23.96 17.84 -23.64 ;
        RECT 15.475 -23.965 15.805 -23.635 ;
        RECT 14.115 -23.965 14.445 -23.635 ;
        RECT 12.755 -23.965 13.085 -23.635 ;
        RECT 11.395 -23.965 11.725 -23.635 ;
        RECT 8.675 -23.965 9.005 -23.635 ;
        RECT 7.315 -23.965 7.645 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -28.04 17.84 -27.72 ;
        RECT 15.475 -28.045 15.805 -27.715 ;
        RECT 14.115 -28.045 14.445 -27.715 ;
        RECT 12.755 -28.045 13.085 -27.715 ;
        RECT 11.395 -28.045 11.725 -27.715 ;
        RECT 8.675 -28.045 9.005 -27.715 ;
        RECT 7.315 -28.045 7.645 -27.715 ;
        RECT 5.955 -28.045 6.285 -27.715 ;
        RECT 4.595 -28.045 4.925 -27.715 ;
        RECT 3.235 -28.045 3.565 -27.715 ;
        RECT 1.875 -28.045 2.205 -27.715 ;
        RECT 0.515 -28.045 0.845 -27.715 ;
        RECT -0.845 -28.045 -0.515 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.72 -34.84 17.84 -34.52 ;
        RECT 16.835 -34.845 17.165 -34.515 ;
        RECT 15.475 -34.845 15.805 -34.515 ;
        RECT 14.115 -34.845 14.445 -34.515 ;
        RECT 12.755 -34.845 13.085 -34.515 ;
        RECT 11.395 -34.845 11.725 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.52 -26.68 21.92 -26.36 ;
        RECT 19.555 -26.685 19.885 -26.355 ;
        RECT 15.475 -26.685 15.805 -26.355 ;
        RECT 14.115 -26.685 14.445 -26.355 ;
        RECT 12.755 -26.685 13.085 -26.355 ;
        RECT 11.395 -26.685 11.725 -26.355 ;
        RECT 8.675 -26.685 9.005 -26.355 ;
        RECT 7.315 -26.685 7.645 -26.355 ;
        RECT 5.955 -26.685 6.285 -26.355 ;
        RECT 4.595 -26.685 4.925 -26.355 ;
        RECT 3.235 -26.685 3.565 -26.355 ;
        RECT 1.875 -26.685 2.205 -26.355 ;
        RECT 0.515 -26.685 0.845 -26.355 ;
        RECT -0.845 -26.685 -0.515 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.68 -29.4 32.12 -29.08 ;
        RECT 30.435 -29.405 30.765 -29.075 ;
        RECT 29.075 -29.405 29.405 -29.075 ;
        RECT 27.715 -29.405 28.045 -29.075 ;
        RECT 26.355 -29.405 26.685 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.6 -23.96 32.8 -23.64 ;
        RECT 30.435 -23.965 30.765 -23.635 ;
        RECT 29.075 -23.965 29.405 -23.635 ;
        RECT 27.715 -23.965 28.045 -23.635 ;
        RECT 26.355 -23.965 26.685 -23.635 ;
        RECT 22.275 -23.965 22.605 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.28 -28.04 32.8 -27.72 ;
        RECT 30.435 -28.045 30.765 -27.715 ;
        RECT 29.075 -28.045 29.405 -27.715 ;
        RECT 27.715 -28.045 28.045 -27.715 ;
        RECT 26.355 -28.045 26.685 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.68 -34.84 32.8 -34.52 ;
        RECT 31.795 -34.845 32.125 -34.515 ;
        RECT 30.435 -34.845 30.765 -34.515 ;
        RECT 29.075 -34.845 29.405 -34.515 ;
        RECT 27.715 -34.845 28.045 -34.515 ;
        RECT 26.355 -34.845 26.685 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.68 -26.68 36.88 -26.36 ;
        RECT 34.515 -26.685 34.845 -26.355 ;
        RECT 30.435 -26.685 30.765 -26.355 ;
        RECT 29.075 -26.685 29.405 -26.355 ;
        RECT 27.715 -26.685 28.045 -26.355 ;
        RECT 26.355 -26.685 26.685 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.64 -29.4 47.08 -29.08 ;
        RECT 45.395 -29.405 45.725 -29.075 ;
        RECT 44.035 -29.405 44.365 -29.075 ;
        RECT 42.675 -29.405 43.005 -29.075 ;
        RECT 41.315 -29.405 41.645 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.56 -23.96 47.76 -23.64 ;
        RECT 45.395 -23.965 45.725 -23.635 ;
        RECT 44.035 -23.965 44.365 -23.635 ;
        RECT 42.675 -23.965 43.005 -23.635 ;
        RECT 41.315 -23.965 41.645 -23.635 ;
        RECT 37.235 -23.965 37.565 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.24 -28.04 47.76 -27.72 ;
        RECT 45.395 -28.045 45.725 -27.715 ;
        RECT 44.035 -28.045 44.365 -27.715 ;
        RECT 42.675 -28.045 43.005 -27.715 ;
        RECT 41.315 -28.045 41.645 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.64 -34.84 47.76 -34.52 ;
        RECT 46.755 -34.845 47.085 -34.515 ;
        RECT 45.395 -34.845 45.725 -34.515 ;
        RECT 44.035 -34.845 44.365 -34.515 ;
        RECT 42.675 -34.845 43.005 -34.515 ;
        RECT 41.315 -34.845 41.645 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.64 -26.68 51.84 -26.36 ;
        RECT 49.475 -26.685 49.805 -26.355 ;
        RECT 45.395 -26.685 45.725 -26.355 ;
        RECT 44.035 -26.685 44.365 -26.355 ;
        RECT 42.675 -26.685 43.005 -26.355 ;
        RECT 41.315 -26.685 41.645 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.6 -29.4 62.04 -29.08 ;
        RECT 60.355 -29.405 60.685 -29.075 ;
        RECT 58.995 -29.405 59.325 -29.075 ;
        RECT 57.635 -29.405 57.965 -29.075 ;
        RECT 56.275 -29.405 56.605 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.52 -23.96 62.72 -23.64 ;
        RECT 60.355 -23.965 60.685 -23.635 ;
        RECT 58.995 -23.965 59.325 -23.635 ;
        RECT 57.635 -23.965 57.965 -23.635 ;
        RECT 56.275 -23.965 56.605 -23.635 ;
        RECT 52.195 -23.965 52.525 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.2 -28.04 62.72 -27.72 ;
        RECT 60.355 -28.045 60.685 -27.715 ;
        RECT 58.995 -28.045 59.325 -27.715 ;
        RECT 57.635 -28.045 57.965 -27.715 ;
        RECT 56.275 -28.045 56.605 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.6 -34.84 62.72 -34.52 ;
        RECT 61.715 -34.845 62.045 -34.515 ;
        RECT 60.355 -34.845 60.685 -34.515 ;
        RECT 58.995 -34.845 59.325 -34.515 ;
        RECT 57.635 -34.845 57.965 -34.515 ;
        RECT 56.275 -34.845 56.605 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.6 -26.68 66.12 -26.36 ;
        RECT 64.435 -26.685 64.765 -26.355 ;
        RECT 60.355 -26.685 60.685 -26.355 ;
        RECT 58.995 -26.685 59.325 -26.355 ;
        RECT 57.635 -26.685 57.965 -26.355 ;
        RECT 56.275 -26.685 56.605 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.56 -29.4 77 -29.08 ;
        RECT 75.315 -29.405 75.645 -29.075 ;
        RECT 73.955 -29.405 74.285 -29.075 ;
        RECT 72.595 -29.405 72.925 -29.075 ;
        RECT 71.235 -29.405 71.565 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.48 -23.96 77.68 -23.64 ;
        RECT 75.315 -23.965 75.645 -23.635 ;
        RECT 73.955 -23.965 74.285 -23.635 ;
        RECT 72.595 -23.965 72.925 -23.635 ;
        RECT 71.235 -23.965 71.565 -23.635 ;
        RECT 67.155 -23.965 67.485 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.16 -28.04 77.68 -27.72 ;
        RECT 75.315 -28.045 75.645 -27.715 ;
        RECT 73.955 -28.045 74.285 -27.715 ;
        RECT 72.595 -28.045 72.925 -27.715 ;
        RECT 71.235 -28.045 71.565 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.56 -34.84 77.68 -34.52 ;
        RECT 76.675 -34.845 77.005 -34.515 ;
        RECT 75.315 -34.845 75.645 -34.515 ;
        RECT 73.955 -34.845 74.285 -34.515 ;
        RECT 72.595 -34.845 72.925 -34.515 ;
        RECT 71.235 -34.845 71.565 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.56 -26.68 81.08 -26.36 ;
        RECT 79.395 -26.685 79.725 -26.355 ;
        RECT 75.315 -26.685 75.645 -26.355 ;
        RECT 73.955 -26.685 74.285 -26.355 ;
        RECT 72.595 -26.685 72.925 -26.355 ;
        RECT 71.235 -26.685 71.565 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.52 -29.4 91.96 -29.08 ;
        RECT 90.275 -29.405 90.605 -29.075 ;
        RECT 88.915 -29.405 89.245 -29.075 ;
        RECT 87.555 -29.405 87.885 -29.075 ;
        RECT 86.195 -29.405 86.525 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.44 -23.96 92.64 -23.64 ;
        RECT 90.275 -23.965 90.605 -23.635 ;
        RECT 88.915 -23.965 89.245 -23.635 ;
        RECT 87.555 -23.965 87.885 -23.635 ;
        RECT 86.195 -23.965 86.525 -23.635 ;
        RECT 82.115 -23.965 82.445 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.12 -28.04 92.64 -27.72 ;
        RECT 90.275 -28.045 90.605 -27.715 ;
        RECT 88.915 -28.045 89.245 -27.715 ;
        RECT 87.555 -28.045 87.885 -27.715 ;
        RECT 86.195 -28.045 86.525 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.52 -34.84 92.64 -34.52 ;
        RECT 91.635 -34.845 91.965 -34.515 ;
        RECT 90.275 -34.845 90.605 -34.515 ;
        RECT 88.915 -34.845 89.245 -34.515 ;
        RECT 87.555 -34.845 87.885 -34.515 ;
        RECT 86.195 -34.845 86.525 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.52 -26.68 96.04 -26.36 ;
        RECT 94.355 -26.685 94.685 -26.355 ;
        RECT 90.275 -26.685 90.605 -26.355 ;
        RECT 88.915 -26.685 89.245 -26.355 ;
        RECT 87.555 -26.685 87.885 -26.355 ;
        RECT 86.195 -26.685 86.525 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.48 -29.4 106.92 -29.08 ;
        RECT 105.235 -29.405 105.565 -29.075 ;
        RECT 103.875 -29.405 104.205 -29.075 ;
        RECT 102.515 -29.405 102.845 -29.075 ;
        RECT 101.155 -29.405 101.485 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.72 -23.96 107.6 -23.64 ;
        RECT 105.235 -23.965 105.565 -23.635 ;
        RECT 103.875 -23.965 104.205 -23.635 ;
        RECT 102.515 -23.965 102.845 -23.635 ;
        RECT 101.155 -23.965 101.485 -23.635 ;
        RECT 97.075 -23.965 97.405 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.4 -28.04 107.6 -27.72 ;
        RECT 105.235 -28.045 105.565 -27.715 ;
        RECT 103.875 -28.045 104.205 -27.715 ;
        RECT 102.515 -28.045 102.845 -27.715 ;
        RECT 101.155 -28.045 101.485 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.48 -34.84 107.6 -34.52 ;
        RECT 106.595 -34.845 106.925 -34.515 ;
        RECT 105.235 -34.845 105.565 -34.515 ;
        RECT 103.875 -34.845 104.205 -34.515 ;
        RECT 102.515 -34.845 102.845 -34.515 ;
        RECT 101.155 -34.845 101.485 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.48 -26.68 111 -26.36 ;
        RECT 109.315 -26.685 109.645 -26.355 ;
        RECT 105.235 -26.685 105.565 -26.355 ;
        RECT 103.875 -26.685 104.205 -26.355 ;
        RECT 102.515 -26.685 102.845 -26.355 ;
        RECT 101.155 -26.685 101.485 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.44 -29.4 121.88 -29.08 ;
        RECT 120.195 -29.405 120.525 -29.075 ;
        RECT 118.835 -29.405 119.165 -29.075 ;
        RECT 117.475 -29.405 117.805 -29.075 ;
        RECT 116.115 -29.405 116.445 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.68 -23.96 122.56 -23.64 ;
        RECT 120.195 -23.965 120.525 -23.635 ;
        RECT 118.835 -23.965 119.165 -23.635 ;
        RECT 117.475 -23.965 117.805 -23.635 ;
        RECT 116.115 -23.965 116.445 -23.635 ;
        RECT 112.035 -23.965 112.365 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.36 -28.04 122.56 -27.72 ;
        RECT 120.195 -28.045 120.525 -27.715 ;
        RECT 118.835 -28.045 119.165 -27.715 ;
        RECT 117.475 -28.045 117.805 -27.715 ;
        RECT 116.115 -28.045 116.445 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.44 -34.84 122.56 -34.52 ;
        RECT 121.555 -34.845 121.885 -34.515 ;
        RECT 120.195 -34.845 120.525 -34.515 ;
        RECT 118.835 -34.845 119.165 -34.515 ;
        RECT 117.475 -34.845 117.805 -34.515 ;
        RECT 116.115 -34.845 116.445 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.44 -26.68 125.96 -26.36 ;
        RECT 124.275 -26.685 124.605 -26.355 ;
        RECT 120.195 -26.685 120.525 -26.355 ;
        RECT 118.835 -26.685 119.165 -26.355 ;
        RECT 117.475 -26.685 117.805 -26.355 ;
        RECT 116.115 -26.685 116.445 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.64 -23.96 136.84 -23.64 ;
        RECT 135.155 -23.965 135.485 -23.635 ;
        RECT 133.795 -23.965 134.125 -23.635 ;
        RECT 132.435 -23.965 132.765 -23.635 ;
        RECT 131.075 -23.965 131.405 -23.635 ;
        RECT 126.995 -23.965 127.325 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.32 -28.04 136.84 -27.72 ;
        RECT 135.155 -28.045 135.485 -27.715 ;
        RECT 133.795 -28.045 134.125 -27.715 ;
        RECT 132.435 -28.045 132.765 -27.715 ;
        RECT 131.075 -28.045 131.405 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.4 -29.4 136.84 -29.08 ;
        RECT 135.155 -29.405 135.485 -29.075 ;
        RECT 133.795 -29.405 134.125 -29.075 ;
        RECT 132.435 -29.405 132.765 -29.075 ;
        RECT 131.075 -29.405 131.405 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -34.845 136.845 -34.515 ;
        RECT 130.4 -34.84 136.845 -34.52 ;
        RECT 135.155 -34.845 135.485 -34.515 ;
        RECT 133.795 -34.845 134.125 -34.515 ;
        RECT 132.435 -34.845 132.765 -34.515 ;
        RECT 131.075 -34.845 131.405 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.4 -26.68 140.92 -26.36 ;
        RECT 139.235 -26.685 139.565 -26.355 ;
        RECT 135.155 -26.685 135.485 -26.355 ;
        RECT 133.795 -26.685 134.125 -26.355 ;
        RECT 132.435 -26.685 132.765 -26.355 ;
        RECT 131.075 -26.685 131.405 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.36 -29.4 151.12 -29.08 ;
        RECT 150.115 -29.405 150.445 -29.075 ;
        RECT 148.755 -29.405 149.085 -29.075 ;
        RECT 147.395 -29.405 147.725 -29.075 ;
        RECT 146.035 -29.405 146.365 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -23.96 151.8 -23.64 ;
        RECT 150.115 -23.965 150.445 -23.635 ;
        RECT 148.755 -23.965 149.085 -23.635 ;
        RECT 147.395 -23.965 147.725 -23.635 ;
        RECT 146.035 -23.965 146.365 -23.635 ;
        RECT 141.955 -23.965 142.285 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.28 -28.04 151.8 -27.72 ;
        RECT 150.115 -28.045 150.445 -27.715 ;
        RECT 148.755 -28.045 149.085 -27.715 ;
        RECT 147.395 -28.045 147.725 -27.715 ;
        RECT 146.035 -28.045 146.365 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -34.845 151.805 -34.515 ;
        RECT 145.36 -34.84 151.805 -34.52 ;
        RECT 150.115 -34.845 150.445 -34.515 ;
        RECT 148.755 -34.845 149.085 -34.515 ;
        RECT 147.395 -34.845 147.725 -34.515 ;
        RECT 146.035 -34.845 146.365 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.36 -26.68 155.88 -26.36 ;
        RECT 154.195 -26.685 154.525 -26.355 ;
        RECT 152.835 -26.685 153.165 -26.355 ;
        RECT 150.115 -26.685 150.445 -26.355 ;
        RECT 148.755 -26.685 149.085 -26.355 ;
        RECT 147.395 -26.685 147.725 -26.355 ;
        RECT 146.035 -26.685 146.365 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.32 -29.4 166.08 -29.08 ;
        RECT 165.075 -29.405 165.405 -29.075 ;
        RECT 163.715 -29.405 164.045 -29.075 ;
        RECT 162.355 -29.405 162.685 -29.075 ;
        RECT 160.995 -29.405 161.325 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.56 -23.96 166.76 -23.64 ;
        RECT 165.075 -23.965 165.405 -23.635 ;
        RECT 163.715 -23.965 164.045 -23.635 ;
        RECT 162.355 -23.965 162.685 -23.635 ;
        RECT 160.995 -23.965 161.325 -23.635 ;
        RECT 156.915 -23.965 157.245 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.24 -28.04 166.76 -27.72 ;
        RECT 165.075 -28.045 165.405 -27.715 ;
        RECT 163.715 -28.045 164.045 -27.715 ;
        RECT 162.355 -28.045 162.685 -27.715 ;
        RECT 160.995 -28.045 161.325 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -34.845 166.765 -34.515 ;
        RECT 160.32 -34.84 166.765 -34.52 ;
        RECT 165.075 -34.845 165.405 -34.515 ;
        RECT 163.715 -34.845 164.045 -34.515 ;
        RECT 162.355 -34.845 162.685 -34.515 ;
        RECT 160.995 -34.845 161.325 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.32 -26.68 170.84 -26.36 ;
        RECT 169.155 -26.685 169.485 -26.355 ;
        RECT 167.795 -26.685 168.125 -26.355 ;
        RECT 165.075 -26.685 165.405 -26.355 ;
        RECT 163.715 -26.685 164.045 -26.355 ;
        RECT 162.355 -26.685 162.685 -26.355 ;
        RECT 160.995 -26.685 161.325 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.28 -29.4 181.04 -29.08 ;
        RECT 180.035 -29.405 180.365 -29.075 ;
        RECT 178.675 -29.405 179.005 -29.075 ;
        RECT 177.315 -29.405 177.645 -29.075 ;
        RECT 175.955 -29.405 176.285 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.52 -23.96 181.72 -23.64 ;
        RECT 180.035 -23.965 180.365 -23.635 ;
        RECT 178.675 -23.965 179.005 -23.635 ;
        RECT 177.315 -23.965 177.645 -23.635 ;
        RECT 175.955 -23.965 176.285 -23.635 ;
        RECT 171.875 -23.965 172.205 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.2 -28.04 181.72 -27.72 ;
        RECT 180.035 -28.045 180.365 -27.715 ;
        RECT 178.675 -28.045 179.005 -27.715 ;
        RECT 177.315 -28.045 177.645 -27.715 ;
        RECT 175.955 -28.045 176.285 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -34.845 181.725 -34.515 ;
        RECT 175.28 -34.84 181.725 -34.52 ;
        RECT 180.035 -34.845 180.365 -34.515 ;
        RECT 178.675 -34.845 179.005 -34.515 ;
        RECT 177.315 -34.845 177.645 -34.515 ;
        RECT 175.955 -34.845 176.285 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.28 -26.68 185.8 -26.36 ;
        RECT 184.115 -26.685 184.445 -26.355 ;
        RECT 182.755 -26.685 183.085 -26.355 ;
        RECT 180.035 -26.685 180.365 -26.355 ;
        RECT 178.675 -26.685 179.005 -26.355 ;
        RECT 177.315 -26.685 177.645 -26.355 ;
        RECT 175.955 -26.685 176.285 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.56 -29.4 196 -29.08 ;
        RECT 194.995 -29.405 195.325 -29.075 ;
        RECT 193.635 -29.405 193.965 -29.075 ;
        RECT 192.275 -29.405 192.605 -29.075 ;
        RECT 190.915 -29.405 191.245 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.48 -23.96 196.68 -23.64 ;
        RECT 194.995 -23.965 195.325 -23.635 ;
        RECT 193.635 -23.965 193.965 -23.635 ;
        RECT 192.275 -23.965 192.605 -23.635 ;
        RECT 190.915 -23.965 191.245 -23.635 ;
        RECT 189.555 -23.965 189.885 -23.635 ;
        RECT 186.835 -23.965 187.165 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.16 -28.04 196.68 -27.72 ;
        RECT 194.995 -28.045 195.325 -27.715 ;
        RECT 193.635 -28.045 193.965 -27.715 ;
        RECT 192.275 -28.045 192.605 -27.715 ;
        RECT 190.915 -28.045 191.245 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -34.845 196.685 -34.515 ;
        RECT 189.56 -34.84 196.685 -34.52 ;
        RECT 194.995 -34.845 195.325 -34.515 ;
        RECT 193.635 -34.845 193.965 -34.515 ;
        RECT 192.275 -34.845 192.605 -34.515 ;
        RECT 190.915 -34.845 191.245 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.56 -26.68 200.76 -26.36 ;
        RECT 199.075 -26.685 199.405 -26.355 ;
        RECT 197.715 -26.685 198.045 -26.355 ;
        RECT 194.995 -26.685 195.325 -26.355 ;
        RECT 193.635 -26.685 193.965 -26.355 ;
        RECT 192.275 -26.685 192.605 -26.355 ;
        RECT 190.915 -26.685 191.245 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.52 -29.4 210.96 -29.08 ;
        RECT 209.955 -29.405 210.285 -29.075 ;
        RECT 208.595 -29.405 208.925 -29.075 ;
        RECT 207.235 -29.405 207.565 -29.075 ;
        RECT 205.875 -29.405 206.205 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.44 -23.96 211.64 -23.64 ;
        RECT 209.955 -23.965 210.285 -23.635 ;
        RECT 208.595 -23.965 208.925 -23.635 ;
        RECT 207.235 -23.965 207.565 -23.635 ;
        RECT 205.875 -23.965 206.205 -23.635 ;
        RECT 204.515 -23.965 204.845 -23.635 ;
        RECT 201.795 -23.965 202.125 -23.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.12 -28.04 211.64 -27.72 ;
        RECT 209.955 -28.045 210.285 -27.715 ;
        RECT 208.595 -28.045 208.925 -27.715 ;
        RECT 207.235 -28.045 207.565 -27.715 ;
        RECT 205.875 -28.045 206.205 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 -34.845 211.645 -34.515 ;
        RECT 204.52 -34.84 211.645 -34.52 ;
        RECT 209.955 -34.845 210.285 -34.515 ;
        RECT 208.595 -34.845 208.925 -34.515 ;
        RECT 207.235 -34.845 207.565 -34.515 ;
        RECT 205.875 -34.845 206.205 -34.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.52 -26.68 215.72 -26.36 ;
        RECT 214.035 -26.685 214.365 -26.355 ;
        RECT 212.675 -26.685 213.005 -26.355 ;
        RECT 209.955 -26.685 210.285 -26.355 ;
        RECT 208.595 -26.685 208.925 -26.355 ;
        RECT 207.235 -26.685 207.565 -26.355 ;
        RECT 205.875 -26.685 206.205 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 -29.405 222.525 -29.075 ;
        RECT 220.835 -29.405 221.165 -29.075 ;
        RECT 219.48 -29.4 225.92 -29.08 ;
        RECT 224.915 -29.405 225.245 -29.075 ;
        RECT 223.555 -29.405 223.885 -29.075 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 954.555 -32.805 954.885 -32.475 ;
        RECT -1.525 -32.8 954.885 -32.48 ;
        RECT 953.195 -32.805 953.525 -32.475 ;
        RECT 951.835 -32.805 952.165 -32.475 ;
        RECT 950.475 -32.805 950.805 -32.475 ;
        RECT 946.395 -32.805 946.725 -32.475 ;
        RECT 945.035 -32.805 945.365 -32.475 ;
        RECT 943.675 -32.805 944.005 -32.475 ;
        RECT 942.315 -32.805 942.645 -32.475 ;
        RECT 940.955 -32.805 941.285 -32.475 ;
        RECT 939.595 -32.805 939.925 -32.475 ;
        RECT 938.235 -32.805 938.565 -32.475 ;
        RECT 936.875 -32.805 937.205 -32.475 ;
        RECT 935.515 -32.805 935.845 -32.475 ;
        RECT 932.795 -32.805 933.125 -32.475 ;
        RECT 930.075 -32.805 930.405 -32.475 ;
        RECT 927.355 -32.805 927.685 -32.475 ;
        RECT 925.995 -32.805 926.325 -32.475 ;
        RECT 924.635 -32.805 924.965 -32.475 ;
        RECT 923.275 -32.805 923.605 -32.475 ;
        RECT 921.915 -32.805 922.245 -32.475 ;
        RECT 920.555 -32.805 920.885 -32.475 ;
        RECT 917.835 -32.805 918.165 -32.475 ;
        RECT 915.115 -32.805 915.445 -32.475 ;
        RECT 912.395 -32.805 912.725 -32.475 ;
        RECT 911.035 -32.805 911.365 -32.475 ;
        RECT 909.675 -32.805 910.005 -32.475 ;
        RECT 908.315 -32.805 908.645 -32.475 ;
        RECT 906.955 -32.805 907.285 -32.475 ;
        RECT 905.595 -32.805 905.925 -32.475 ;
        RECT 902.875 -32.805 903.205 -32.475 ;
        RECT 900.155 -32.805 900.485 -32.475 ;
        RECT 897.435 -32.805 897.765 -32.475 ;
        RECT 896.075 -32.805 896.405 -32.475 ;
        RECT 894.715 -32.805 895.045 -32.475 ;
        RECT 893.355 -32.805 893.685 -32.475 ;
        RECT 891.995 -32.805 892.325 -32.475 ;
        RECT 890.635 -32.805 890.965 -32.475 ;
        RECT 887.915 -32.805 888.245 -32.475 ;
        RECT 885.195 -32.805 885.525 -32.475 ;
        RECT 882.475 -32.805 882.805 -32.475 ;
        RECT 881.115 -32.805 881.445 -32.475 ;
        RECT 879.755 -32.805 880.085 -32.475 ;
        RECT 878.395 -32.805 878.725 -32.475 ;
        RECT 877.035 -32.805 877.365 -32.475 ;
        RECT 875.675 -32.805 876.005 -32.475 ;
        RECT 872.955 -32.805 873.285 -32.475 ;
        RECT 870.235 -32.805 870.565 -32.475 ;
        RECT 867.515 -32.805 867.845 -32.475 ;
        RECT 866.155 -32.805 866.485 -32.475 ;
        RECT 864.795 -32.805 865.125 -32.475 ;
        RECT 863.435 -32.805 863.765 -32.475 ;
        RECT 862.075 -32.805 862.405 -32.475 ;
        RECT 860.715 -32.805 861.045 -32.475 ;
        RECT 857.995 -32.805 858.325 -32.475 ;
        RECT 855.275 -32.805 855.605 -32.475 ;
        RECT 852.555 -32.805 852.885 -32.475 ;
        RECT 851.195 -32.805 851.525 -32.475 ;
        RECT 849.835 -32.805 850.165 -32.475 ;
        RECT 848.475 -32.805 848.805 -32.475 ;
        RECT 847.115 -32.805 847.445 -32.475 ;
        RECT 845.755 -32.805 846.085 -32.475 ;
        RECT 843.035 -32.805 843.365 -32.475 ;
        RECT 840.315 -32.805 840.645 -32.475 ;
        RECT 837.595 -32.805 837.925 -32.475 ;
        RECT 836.235 -32.805 836.565 -32.475 ;
        RECT 834.875 -32.805 835.205 -32.475 ;
        RECT 833.515 -32.805 833.845 -32.475 ;
        RECT 832.155 -32.805 832.485 -32.475 ;
        RECT 828.075 -32.805 828.405 -32.475 ;
        RECT 825.355 -32.805 825.685 -32.475 ;
        RECT 822.635 -32.805 822.965 -32.475 ;
        RECT 821.275 -32.805 821.605 -32.475 ;
        RECT 819.915 -32.805 820.245 -32.475 ;
        RECT 818.555 -32.805 818.885 -32.475 ;
        RECT 817.195 -32.805 817.525 -32.475 ;
        RECT 813.115 -32.805 813.445 -32.475 ;
        RECT 810.395 -32.805 810.725 -32.475 ;
        RECT 807.675 -32.805 808.005 -32.475 ;
        RECT 806.315 -32.805 806.645 -32.475 ;
        RECT 804.955 -32.805 805.285 -32.475 ;
        RECT 803.595 -32.805 803.925 -32.475 ;
        RECT 802.235 -32.805 802.565 -32.475 ;
        RECT 798.155 -32.805 798.485 -32.475 ;
        RECT 795.435 -32.805 795.765 -32.475 ;
        RECT 792.715 -32.805 793.045 -32.475 ;
        RECT 791.355 -32.805 791.685 -32.475 ;
        RECT 789.995 -32.805 790.325 -32.475 ;
        RECT 788.635 -32.805 788.965 -32.475 ;
        RECT 787.275 -32.805 787.605 -32.475 ;
        RECT 783.195 -32.805 783.525 -32.475 ;
        RECT 780.475 -32.805 780.805 -32.475 ;
        RECT 779.115 -32.805 779.445 -32.475 ;
        RECT 777.755 -32.805 778.085 -32.475 ;
        RECT 776.395 -32.805 776.725 -32.475 ;
        RECT 775.035 -32.805 775.365 -32.475 ;
        RECT 773.675 -32.805 774.005 -32.475 ;
        RECT 772.315 -32.805 772.645 -32.475 ;
        RECT 768.235 -32.805 768.565 -32.475 ;
        RECT 764.155 -32.805 764.485 -32.475 ;
        RECT 762.795 -32.805 763.125 -32.475 ;
        RECT 761.435 -32.805 761.765 -32.475 ;
        RECT 760.075 -32.805 760.405 -32.475 ;
        RECT 758.715 -32.805 759.045 -32.475 ;
        RECT 757.355 -32.805 757.685 -32.475 ;
        RECT 753.275 -32.805 753.605 -32.475 ;
        RECT 749.195 -32.805 749.525 -32.475 ;
        RECT 747.835 -32.805 748.165 -32.475 ;
        RECT 746.475 -32.805 746.805 -32.475 ;
        RECT 745.115 -32.805 745.445 -32.475 ;
        RECT 743.755 -32.805 744.085 -32.475 ;
        RECT 742.395 -32.805 742.725 -32.475 ;
        RECT 738.315 -32.805 738.645 -32.475 ;
        RECT 734.235 -32.805 734.565 -32.475 ;
        RECT 732.875 -32.805 733.205 -32.475 ;
        RECT 731.515 -32.805 731.845 -32.475 ;
        RECT 730.155 -32.805 730.485 -32.475 ;
        RECT 728.795 -32.805 729.125 -32.475 ;
        RECT 727.435 -32.805 727.765 -32.475 ;
        RECT 721.995 -32.805 722.325 -32.475 ;
        RECT 719.275 -32.805 719.605 -32.475 ;
        RECT 717.915 -32.805 718.245 -32.475 ;
        RECT 716.555 -32.805 716.885 -32.475 ;
        RECT 715.195 -32.805 715.525 -32.475 ;
        RECT 713.835 -32.805 714.165 -32.475 ;
        RECT 712.475 -32.805 712.805 -32.475 ;
        RECT 707.035 -32.805 707.365 -32.475 ;
        RECT 704.315 -32.805 704.645 -32.475 ;
        RECT 702.955 -32.805 703.285 -32.475 ;
        RECT 701.595 -32.805 701.925 -32.475 ;
        RECT 700.235 -32.805 700.565 -32.475 ;
        RECT 698.875 -32.805 699.205 -32.475 ;
        RECT 697.515 -32.805 697.845 -32.475 ;
        RECT 692.075 -32.805 692.405 -32.475 ;
        RECT 689.355 -32.805 689.685 -32.475 ;
        RECT 687.995 -32.805 688.325 -32.475 ;
        RECT 686.635 -32.805 686.965 -32.475 ;
        RECT 685.275 -32.805 685.605 -32.475 ;
        RECT 683.915 -32.805 684.245 -32.475 ;
        RECT 682.555 -32.805 682.885 -32.475 ;
        RECT 679.835 -32.805 680.165 -32.475 ;
        RECT 677.115 -32.805 677.445 -32.475 ;
        RECT 674.395 -32.805 674.725 -32.475 ;
        RECT 673.035 -32.805 673.365 -32.475 ;
        RECT 671.675 -32.805 672.005 -32.475 ;
        RECT 670.315 -32.805 670.645 -32.475 ;
        RECT 668.955 -32.805 669.285 -32.475 ;
        RECT 667.595 -32.805 667.925 -32.475 ;
        RECT 664.875 -32.805 665.205 -32.475 ;
        RECT 662.155 -32.805 662.485 -32.475 ;
        RECT 659.435 -32.805 659.765 -32.475 ;
        RECT 658.075 -32.805 658.405 -32.475 ;
        RECT 656.715 -32.805 657.045 -32.475 ;
        RECT 655.355 -32.805 655.685 -32.475 ;
        RECT 653.995 -32.805 654.325 -32.475 ;
        RECT 652.635 -32.805 652.965 -32.475 ;
        RECT 649.915 -32.805 650.245 -32.475 ;
        RECT 647.195 -32.805 647.525 -32.475 ;
        RECT 644.475 -32.805 644.805 -32.475 ;
        RECT 643.115 -32.805 643.445 -32.475 ;
        RECT 641.755 -32.805 642.085 -32.475 ;
        RECT 640.395 -32.805 640.725 -32.475 ;
        RECT 639.035 -32.805 639.365 -32.475 ;
        RECT 637.675 -32.805 638.005 -32.475 ;
        RECT 634.955 -32.805 635.285 -32.475 ;
        RECT 632.235 -32.805 632.565 -32.475 ;
        RECT 629.515 -32.805 629.845 -32.475 ;
        RECT 628.155 -32.805 628.485 -32.475 ;
        RECT 626.795 -32.805 627.125 -32.475 ;
        RECT 625.435 -32.805 625.765 -32.475 ;
        RECT 624.075 -32.805 624.405 -32.475 ;
        RECT 622.715 -32.805 623.045 -32.475 ;
        RECT 619.995 -32.805 620.325 -32.475 ;
        RECT 617.275 -32.805 617.605 -32.475 ;
        RECT 614.555 -32.805 614.885 -32.475 ;
        RECT 613.195 -32.805 613.525 -32.475 ;
        RECT 611.835 -32.805 612.165 -32.475 ;
        RECT 610.475 -32.805 610.805 -32.475 ;
        RECT 609.115 -32.805 609.445 -32.475 ;
        RECT 607.755 -32.805 608.085 -32.475 ;
        RECT 605.035 -32.805 605.365 -32.475 ;
        RECT 602.315 -32.805 602.645 -32.475 ;
        RECT 599.595 -32.805 599.925 -32.475 ;
        RECT 598.235 -32.805 598.565 -32.475 ;
        RECT 596.875 -32.805 597.205 -32.475 ;
        RECT 595.515 -32.805 595.845 -32.475 ;
        RECT 594.155 -32.805 594.485 -32.475 ;
        RECT 592.795 -32.805 593.125 -32.475 ;
        RECT 590.075 -32.805 590.405 -32.475 ;
        RECT 587.355 -32.805 587.685 -32.475 ;
        RECT 584.635 -32.805 584.965 -32.475 ;
        RECT 583.275 -32.805 583.605 -32.475 ;
        RECT 581.915 -32.805 582.245 -32.475 ;
        RECT 580.555 -32.805 580.885 -32.475 ;
        RECT 579.195 -32.805 579.525 -32.475 ;
        RECT 577.835 -32.805 578.165 -32.475 ;
        RECT 575.115 -32.805 575.445 -32.475 ;
        RECT 572.395 -32.805 572.725 -32.475 ;
        RECT 569.675 -32.805 570.005 -32.475 ;
        RECT 568.315 -32.805 568.645 -32.475 ;
        RECT 566.955 -32.805 567.285 -32.475 ;
        RECT 565.595 -32.805 565.925 -32.475 ;
        RECT 564.235 -32.805 564.565 -32.475 ;
        RECT 562.875 -32.805 563.205 -32.475 ;
        RECT 560.155 -32.805 560.485 -32.475 ;
        RECT 557.435 -32.805 557.765 -32.475 ;
        RECT 554.715 -32.805 555.045 -32.475 ;
        RECT 553.355 -32.805 553.685 -32.475 ;
        RECT 551.995 -32.805 552.325 -32.475 ;
        RECT 550.635 -32.805 550.965 -32.475 ;
        RECT 549.275 -32.805 549.605 -32.475 ;
        RECT 547.915 -32.805 548.245 -32.475 ;
        RECT 545.195 -32.805 545.525 -32.475 ;
        RECT 542.475 -32.805 542.805 -32.475 ;
        RECT 539.755 -32.805 540.085 -32.475 ;
        RECT 538.395 -32.805 538.725 -32.475 ;
        RECT 537.035 -32.805 537.365 -32.475 ;
        RECT 535.675 -32.805 536.005 -32.475 ;
        RECT 534.315 -32.805 534.645 -32.475 ;
        RECT 532.955 -32.805 533.285 -32.475 ;
        RECT 530.235 -32.805 530.565 -32.475 ;
        RECT 527.515 -32.805 527.845 -32.475 ;
        RECT 524.795 -32.805 525.125 -32.475 ;
        RECT 523.435 -32.805 523.765 -32.475 ;
        RECT 522.075 -32.805 522.405 -32.475 ;
        RECT 520.715 -32.805 521.045 -32.475 ;
        RECT 519.355 -32.805 519.685 -32.475 ;
        RECT 517.995 -32.805 518.325 -32.475 ;
        RECT 515.275 -32.805 515.605 -32.475 ;
        RECT 512.555 -32.805 512.885 -32.475 ;
        RECT 509.835 -32.805 510.165 -32.475 ;
        RECT 508.475 -32.805 508.805 -32.475 ;
        RECT 507.115 -32.805 507.445 -32.475 ;
        RECT 505.755 -32.805 506.085 -32.475 ;
        RECT 504.395 -32.805 504.725 -32.475 ;
        RECT 500.315 -32.805 500.645 -32.475 ;
        RECT 497.595 -32.805 497.925 -32.475 ;
        RECT 494.875 -32.805 495.205 -32.475 ;
        RECT 493.515 -32.805 493.845 -32.475 ;
        RECT 492.155 -32.805 492.485 -32.475 ;
        RECT 490.795 -32.805 491.125 -32.475 ;
        RECT 489.435 -32.805 489.765 -32.475 ;
        RECT 485.355 -32.805 485.685 -32.475 ;
        RECT 482.635 -32.805 482.965 -32.475 ;
        RECT 479.915 -32.805 480.245 -32.475 ;
        RECT 478.555 -32.805 478.885 -32.475 ;
        RECT 477.195 -32.805 477.525 -32.475 ;
        RECT 475.835 -32.805 476.165 -32.475 ;
        RECT 474.475 -32.805 474.805 -32.475 ;
        RECT 470.395 -32.805 470.725 -32.475 ;
        RECT 467.675 -32.805 468.005 -32.475 ;
        RECT 464.955 -32.805 465.285 -32.475 ;
        RECT 463.595 -32.805 463.925 -32.475 ;
        RECT 462.235 -32.805 462.565 -32.475 ;
        RECT 460.875 -32.805 461.205 -32.475 ;
        RECT 459.515 -32.805 459.845 -32.475 ;
        RECT 455.435 -32.805 455.765 -32.475 ;
        RECT 452.715 -32.805 453.045 -32.475 ;
        RECT 449.995 -32.805 450.325 -32.475 ;
        RECT 448.635 -32.805 448.965 -32.475 ;
        RECT 447.275 -32.805 447.605 -32.475 ;
        RECT 445.915 -32.805 446.245 -32.475 ;
        RECT 444.555 -32.805 444.885 -32.475 ;
        RECT 440.475 -32.805 440.805 -32.475 ;
        RECT 436.395 -32.805 436.725 -32.475 ;
        RECT 435.035 -32.805 435.365 -32.475 ;
        RECT 433.675 -32.805 434.005 -32.475 ;
        RECT 432.315 -32.805 432.645 -32.475 ;
        RECT 430.955 -32.805 431.285 -32.475 ;
        RECT 429.595 -32.805 429.925 -32.475 ;
        RECT 425.515 -32.805 425.845 -32.475 ;
        RECT 421.435 -32.805 421.765 -32.475 ;
        RECT 420.075 -32.805 420.405 -32.475 ;
        RECT 418.715 -32.805 419.045 -32.475 ;
        RECT 417.355 -32.805 417.685 -32.475 ;
        RECT 415.995 -32.805 416.325 -32.475 ;
        RECT 414.635 -32.805 414.965 -32.475 ;
        RECT 410.555 -32.805 410.885 -32.475 ;
        RECT 406.475 -32.805 406.805 -32.475 ;
        RECT 405.115 -32.805 405.445 -32.475 ;
        RECT 403.755 -32.805 404.085 -32.475 ;
        RECT 402.395 -32.805 402.725 -32.475 ;
        RECT 401.035 -32.805 401.365 -32.475 ;
        RECT 399.675 -32.805 400.005 -32.475 ;
        RECT 395.595 -32.805 395.925 -32.475 ;
        RECT 394.235 -32.805 394.565 -32.475 ;
        RECT 391.515 -32.805 391.845 -32.475 ;
        RECT 390.155 -32.805 390.485 -32.475 ;
        RECT 388.795 -32.805 389.125 -32.475 ;
        RECT 387.435 -32.805 387.765 -32.475 ;
        RECT 386.075 -32.805 386.405 -32.475 ;
        RECT 384.715 -32.805 385.045 -32.475 ;
        RECT 379.275 -32.805 379.605 -32.475 ;
        RECT 376.555 -32.805 376.885 -32.475 ;
        RECT 375.195 -32.805 375.525 -32.475 ;
        RECT 373.835 -32.805 374.165 -32.475 ;
        RECT 372.475 -32.805 372.805 -32.475 ;
        RECT 371.115 -32.805 371.445 -32.475 ;
        RECT 369.755 -32.805 370.085 -32.475 ;
        RECT 364.315 -32.805 364.645 -32.475 ;
        RECT 361.595 -32.805 361.925 -32.475 ;
        RECT 360.235 -32.805 360.565 -32.475 ;
        RECT 358.875 -32.805 359.205 -32.475 ;
        RECT 357.515 -32.805 357.845 -32.475 ;
        RECT 356.155 -32.805 356.485 -32.475 ;
        RECT 354.795 -32.805 355.125 -32.475 ;
        RECT 349.355 -32.805 349.685 -32.475 ;
        RECT 346.635 -32.805 346.965 -32.475 ;
        RECT 345.275 -32.805 345.605 -32.475 ;
        RECT 343.915 -32.805 344.245 -32.475 ;
        RECT 342.555 -32.805 342.885 -32.475 ;
        RECT 341.195 -32.805 341.525 -32.475 ;
        RECT 339.835 -32.805 340.165 -32.475 ;
        RECT 337.115 -32.805 337.445 -32.475 ;
        RECT 334.395 -32.805 334.725 -32.475 ;
        RECT 331.675 -32.805 332.005 -32.475 ;
        RECT 330.315 -32.805 330.645 -32.475 ;
        RECT 328.955 -32.805 329.285 -32.475 ;
        RECT 327.595 -32.805 327.925 -32.475 ;
        RECT 326.235 -32.805 326.565 -32.475 ;
        RECT 324.875 -32.805 325.205 -32.475 ;
        RECT 322.155 -32.805 322.485 -32.475 ;
        RECT 319.435 -32.805 319.765 -32.475 ;
        RECT 316.715 -32.805 317.045 -32.475 ;
        RECT 315.355 -32.805 315.685 -32.475 ;
        RECT 313.995 -32.805 314.325 -32.475 ;
        RECT 312.635 -32.805 312.965 -32.475 ;
        RECT 311.275 -32.805 311.605 -32.475 ;
        RECT 309.915 -32.805 310.245 -32.475 ;
        RECT 307.195 -32.805 307.525 -32.475 ;
        RECT 304.475 -32.805 304.805 -32.475 ;
        RECT 301.755 -32.805 302.085 -32.475 ;
        RECT 300.395 -32.805 300.725 -32.475 ;
        RECT 299.035 -32.805 299.365 -32.475 ;
        RECT 297.675 -32.805 298.005 -32.475 ;
        RECT 296.315 -32.805 296.645 -32.475 ;
        RECT 294.955 -32.805 295.285 -32.475 ;
        RECT 292.235 -32.805 292.565 -32.475 ;
        RECT 289.515 -32.805 289.845 -32.475 ;
        RECT 286.795 -32.805 287.125 -32.475 ;
        RECT 285.435 -32.805 285.765 -32.475 ;
        RECT 284.075 -32.805 284.405 -32.475 ;
        RECT 282.715 -32.805 283.045 -32.475 ;
        RECT 281.355 -32.805 281.685 -32.475 ;
        RECT 279.995 -32.805 280.325 -32.475 ;
        RECT 277.275 -32.805 277.605 -32.475 ;
        RECT 274.555 -32.805 274.885 -32.475 ;
        RECT 271.835 -32.805 272.165 -32.475 ;
        RECT 270.475 -32.805 270.805 -32.475 ;
        RECT 269.115 -32.805 269.445 -32.475 ;
        RECT 267.755 -32.805 268.085 -32.475 ;
        RECT 266.395 -32.805 266.725 -32.475 ;
        RECT 265.035 -32.805 265.365 -32.475 ;
        RECT 262.315 -32.805 262.645 -32.475 ;
        RECT 259.595 -32.805 259.925 -32.475 ;
        RECT 256.875 -32.805 257.205 -32.475 ;
        RECT 255.515 -32.805 255.845 -32.475 ;
        RECT 254.155 -32.805 254.485 -32.475 ;
        RECT 252.795 -32.805 253.125 -32.475 ;
        RECT 251.435 -32.805 251.765 -32.475 ;
        RECT 250.075 -32.805 250.405 -32.475 ;
        RECT 247.355 -32.805 247.685 -32.475 ;
        RECT 244.635 -32.805 244.965 -32.475 ;
        RECT 241.915 -32.805 242.245 -32.475 ;
        RECT 240.555 -32.805 240.885 -32.475 ;
        RECT 239.195 -32.805 239.525 -32.475 ;
        RECT 237.835 -32.805 238.165 -32.475 ;
        RECT 236.475 -32.805 236.805 -32.475 ;
        RECT 235.115 -32.805 235.445 -32.475 ;
        RECT 232.395 -32.805 232.725 -32.475 ;
        RECT 229.675 -32.805 230.005 -32.475 ;
        RECT 226.955 -32.805 227.285 -32.475 ;
        RECT 225.595 -32.805 225.925 -32.475 ;
        RECT 224.235 -32.805 224.565 -32.475 ;
        RECT 222.875 -32.805 223.205 -32.475 ;
        RECT 221.515 -32.805 221.845 -32.475 ;
        RECT 220.155 -32.805 220.485 -32.475 ;
        RECT 217.435 -32.805 217.765 -32.475 ;
        RECT 214.715 -32.805 215.045 -32.475 ;
        RECT 211.995 -32.805 212.325 -32.475 ;
        RECT 210.635 -32.805 210.965 -32.475 ;
        RECT 209.275 -32.805 209.605 -32.475 ;
        RECT 207.915 -32.805 208.245 -32.475 ;
        RECT 206.555 -32.805 206.885 -32.475 ;
        RECT 205.195 -32.805 205.525 -32.475 ;
        RECT 202.475 -32.805 202.805 -32.475 ;
        RECT 199.755 -32.805 200.085 -32.475 ;
        RECT 197.035 -32.805 197.365 -32.475 ;
        RECT 195.675 -32.805 196.005 -32.475 ;
        RECT 194.315 -32.805 194.645 -32.475 ;
        RECT 192.955 -32.805 193.285 -32.475 ;
        RECT 191.595 -32.805 191.925 -32.475 ;
        RECT 190.235 -32.805 190.565 -32.475 ;
        RECT 187.515 -32.805 187.845 -32.475 ;
        RECT 184.795 -32.805 185.125 -32.475 ;
        RECT 182.075 -32.805 182.405 -32.475 ;
        RECT 180.715 -32.805 181.045 -32.475 ;
        RECT 179.355 -32.805 179.685 -32.475 ;
        RECT 177.995 -32.805 178.325 -32.475 ;
        RECT 176.635 -32.805 176.965 -32.475 ;
        RECT 175.275 -32.805 175.605 -32.475 ;
        RECT 172.555 -32.805 172.885 -32.475 ;
        RECT 169.835 -32.805 170.165 -32.475 ;
        RECT 167.115 -32.805 167.445 -32.475 ;
        RECT 165.755 -32.805 166.085 -32.475 ;
        RECT 164.395 -32.805 164.725 -32.475 ;
        RECT 163.035 -32.805 163.365 -32.475 ;
        RECT 161.675 -32.805 162.005 -32.475 ;
        RECT 157.595 -32.805 157.925 -32.475 ;
        RECT 154.875 -32.805 155.205 -32.475 ;
        RECT 152.155 -32.805 152.485 -32.475 ;
        RECT 150.795 -32.805 151.125 -32.475 ;
        RECT 149.435 -32.805 149.765 -32.475 ;
        RECT 148.075 -32.805 148.405 -32.475 ;
        RECT 146.715 -32.805 147.045 -32.475 ;
        RECT 142.635 -32.805 142.965 -32.475 ;
        RECT 139.915 -32.805 140.245 -32.475 ;
        RECT 137.195 -32.805 137.525 -32.475 ;
        RECT 135.835 -32.805 136.165 -32.475 ;
        RECT 134.475 -32.805 134.805 -32.475 ;
        RECT 133.115 -32.805 133.445 -32.475 ;
        RECT 131.755 -32.805 132.085 -32.475 ;
        RECT 127.675 -32.805 128.005 -32.475 ;
        RECT 124.955 -32.805 125.285 -32.475 ;
        RECT 122.235 -32.805 122.565 -32.475 ;
        RECT 120.875 -32.805 121.205 -32.475 ;
        RECT 119.515 -32.805 119.845 -32.475 ;
        RECT 118.155 -32.805 118.485 -32.475 ;
        RECT 116.795 -32.805 117.125 -32.475 ;
        RECT 112.715 -32.805 113.045 -32.475 ;
        RECT 109.995 -32.805 110.325 -32.475 ;
        RECT 107.275 -32.805 107.605 -32.475 ;
        RECT 105.915 -32.805 106.245 -32.475 ;
        RECT 104.555 -32.805 104.885 -32.475 ;
        RECT 103.195 -32.805 103.525 -32.475 ;
        RECT 101.835 -32.805 102.165 -32.475 ;
        RECT 97.755 -32.805 98.085 -32.475 ;
        RECT 93.675 -32.805 94.005 -32.475 ;
        RECT 92.315 -32.805 92.645 -32.475 ;
        RECT 90.955 -32.805 91.285 -32.475 ;
        RECT 89.595 -32.805 89.925 -32.475 ;
        RECT 88.235 -32.805 88.565 -32.475 ;
        RECT 86.875 -32.805 87.205 -32.475 ;
        RECT 82.795 -32.805 83.125 -32.475 ;
        RECT 78.715 -32.805 79.045 -32.475 ;
        RECT 77.355 -32.805 77.685 -32.475 ;
        RECT 75.995 -32.805 76.325 -32.475 ;
        RECT 74.635 -32.805 74.965 -32.475 ;
        RECT 73.275 -32.805 73.605 -32.475 ;
        RECT 71.915 -32.805 72.245 -32.475 ;
        RECT 67.835 -32.805 68.165 -32.475 ;
        RECT 63.755 -32.805 64.085 -32.475 ;
        RECT 62.395 -32.805 62.725 -32.475 ;
        RECT 61.035 -32.805 61.365 -32.475 ;
        RECT 59.675 -32.805 60.005 -32.475 ;
        RECT 58.315 -32.805 58.645 -32.475 ;
        RECT 56.955 -32.805 57.285 -32.475 ;
        RECT 51.515 -32.805 51.845 -32.475 ;
        RECT 48.795 -32.805 49.125 -32.475 ;
        RECT 47.435 -32.805 47.765 -32.475 ;
        RECT 46.075 -32.805 46.405 -32.475 ;
        RECT 44.715 -32.805 45.045 -32.475 ;
        RECT 43.355 -32.805 43.685 -32.475 ;
        RECT 41.995 -32.805 42.325 -32.475 ;
        RECT 36.555 -32.805 36.885 -32.475 ;
        RECT 33.835 -32.805 34.165 -32.475 ;
        RECT 32.475 -32.805 32.805 -32.475 ;
        RECT 31.115 -32.805 31.445 -32.475 ;
        RECT 29.755 -32.805 30.085 -32.475 ;
        RECT 28.395 -32.805 28.725 -32.475 ;
        RECT 27.035 -32.805 27.365 -32.475 ;
        RECT 21.595 -32.805 21.925 -32.475 ;
        RECT 18.875 -32.805 19.205 -32.475 ;
        RECT 17.515 -32.805 17.845 -32.475 ;
        RECT 16.155 -32.805 16.485 -32.475 ;
        RECT 14.795 -32.805 15.125 -32.475 ;
        RECT 13.435 -32.805 13.765 -32.475 ;
        RECT 12.075 -32.805 12.405 -32.475 ;
        RECT 10.715 -32.805 11.045 -32.475 ;
        RECT 7.995 -32.805 8.325 -32.475 ;
        RECT 6.635 -32.805 6.965 -32.475 ;
        RECT 5.275 -32.805 5.605 -32.475 ;
        RECT 3.915 -32.805 4.245 -32.475 ;
        RECT 2.555 -32.805 2.885 -32.475 ;
        RECT 1.195 -32.805 1.525 -32.475 ;
        RECT -0.165 -32.805 0.165 -32.475 ;
        RECT -1.525 -32.805 -1.195 -32.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -34.165 954.885 -33.835 ;
        RECT -1.525 -34.16 954.885 -33.84 ;
        RECT 953.195 -34.165 953.525 -33.835 ;
        RECT 951.835 -34.165 952.165 -33.835 ;
        RECT 950.475 -34.165 950.805 -33.835 ;
        RECT 946.395 -34.165 946.725 -33.835 ;
        RECT 945.035 -34.165 945.365 -33.835 ;
        RECT 943.675 -34.165 944.005 -33.835 ;
        RECT 942.315 -34.165 942.645 -33.835 ;
        RECT 940.955 -34.165 941.285 -33.835 ;
        RECT 939.595 -34.165 939.925 -33.835 ;
        RECT 938.235 -34.165 938.565 -33.835 ;
        RECT 936.875 -34.165 937.205 -33.835 ;
        RECT 935.515 -34.165 935.845 -33.835 ;
        RECT 932.795 -34.165 933.125 -33.835 ;
        RECT 930.075 -34.165 930.405 -33.835 ;
        RECT 927.355 -34.165 927.685 -33.835 ;
        RECT 925.995 -34.165 926.325 -33.835 ;
        RECT 924.635 -34.165 924.965 -33.835 ;
        RECT 923.275 -34.165 923.605 -33.835 ;
        RECT 921.915 -34.165 922.245 -33.835 ;
        RECT 920.555 -34.165 920.885 -33.835 ;
        RECT 917.835 -34.165 918.165 -33.835 ;
        RECT 915.115 -34.165 915.445 -33.835 ;
        RECT 912.395 -34.165 912.725 -33.835 ;
        RECT 911.035 -34.165 911.365 -33.835 ;
        RECT 909.675 -34.165 910.005 -33.835 ;
        RECT 908.315 -34.165 908.645 -33.835 ;
        RECT 906.955 -34.165 907.285 -33.835 ;
        RECT 905.595 -34.165 905.925 -33.835 ;
        RECT 902.875 -34.165 903.205 -33.835 ;
        RECT 900.155 -34.165 900.485 -33.835 ;
        RECT 897.435 -34.165 897.765 -33.835 ;
        RECT 896.075 -34.165 896.405 -33.835 ;
        RECT 894.715 -34.165 895.045 -33.835 ;
        RECT 893.355 -34.165 893.685 -33.835 ;
        RECT 891.995 -34.165 892.325 -33.835 ;
        RECT 890.635 -34.165 890.965 -33.835 ;
        RECT 887.915 -34.165 888.245 -33.835 ;
        RECT 885.195 -34.165 885.525 -33.835 ;
        RECT 882.475 -34.165 882.805 -33.835 ;
        RECT 881.115 -34.165 881.445 -33.835 ;
        RECT 879.755 -34.165 880.085 -33.835 ;
        RECT 878.395 -34.165 878.725 -33.835 ;
        RECT 877.035 -34.165 877.365 -33.835 ;
        RECT 875.675 -34.165 876.005 -33.835 ;
        RECT 872.955 -34.165 873.285 -33.835 ;
        RECT 870.235 -34.165 870.565 -33.835 ;
        RECT 867.515 -34.165 867.845 -33.835 ;
        RECT 866.155 -34.165 866.485 -33.835 ;
        RECT 864.795 -34.165 865.125 -33.835 ;
        RECT 863.435 -34.165 863.765 -33.835 ;
        RECT 862.075 -34.165 862.405 -33.835 ;
        RECT 860.715 -34.165 861.045 -33.835 ;
        RECT 857.995 -34.165 858.325 -33.835 ;
        RECT 855.275 -34.165 855.605 -33.835 ;
        RECT 852.555 -34.165 852.885 -33.835 ;
        RECT 851.195 -34.165 851.525 -33.835 ;
        RECT 849.835 -34.165 850.165 -33.835 ;
        RECT 848.475 -34.165 848.805 -33.835 ;
        RECT 847.115 -34.165 847.445 -33.835 ;
        RECT 845.755 -34.165 846.085 -33.835 ;
        RECT 843.035 -34.165 843.365 -33.835 ;
        RECT 840.315 -34.165 840.645 -33.835 ;
        RECT 837.595 -34.165 837.925 -33.835 ;
        RECT 836.235 -34.165 836.565 -33.835 ;
        RECT 834.875 -34.165 835.205 -33.835 ;
        RECT 833.515 -34.165 833.845 -33.835 ;
        RECT 832.155 -34.165 832.485 -33.835 ;
        RECT 828.075 -34.165 828.405 -33.835 ;
        RECT 825.355 -34.165 825.685 -33.835 ;
        RECT 822.635 -34.165 822.965 -33.835 ;
        RECT 821.275 -34.165 821.605 -33.835 ;
        RECT 819.915 -34.165 820.245 -33.835 ;
        RECT 818.555 -34.165 818.885 -33.835 ;
        RECT 817.195 -34.165 817.525 -33.835 ;
        RECT 813.115 -34.165 813.445 -33.835 ;
        RECT 810.395 -34.165 810.725 -33.835 ;
        RECT 807.675 -34.165 808.005 -33.835 ;
        RECT 806.315 -34.165 806.645 -33.835 ;
        RECT 804.955 -34.165 805.285 -33.835 ;
        RECT 803.595 -34.165 803.925 -33.835 ;
        RECT 802.235 -34.165 802.565 -33.835 ;
        RECT 798.155 -34.165 798.485 -33.835 ;
        RECT 795.435 -34.165 795.765 -33.835 ;
        RECT 792.715 -34.165 793.045 -33.835 ;
        RECT 791.355 -34.165 791.685 -33.835 ;
        RECT 789.995 -34.165 790.325 -33.835 ;
        RECT 788.635 -34.165 788.965 -33.835 ;
        RECT 787.275 -34.165 787.605 -33.835 ;
        RECT 783.195 -34.165 783.525 -33.835 ;
        RECT 780.475 -34.165 780.805 -33.835 ;
        RECT 779.115 -34.165 779.445 -33.835 ;
        RECT 777.755 -34.165 778.085 -33.835 ;
        RECT 776.395 -34.165 776.725 -33.835 ;
        RECT 775.035 -34.165 775.365 -33.835 ;
        RECT 773.675 -34.165 774.005 -33.835 ;
        RECT 772.315 -34.165 772.645 -33.835 ;
        RECT 768.235 -34.165 768.565 -33.835 ;
        RECT 764.155 -34.165 764.485 -33.835 ;
        RECT 762.795 -34.165 763.125 -33.835 ;
        RECT 761.435 -34.165 761.765 -33.835 ;
        RECT 760.075 -34.165 760.405 -33.835 ;
        RECT 758.715 -34.165 759.045 -33.835 ;
        RECT 757.355 -34.165 757.685 -33.835 ;
        RECT 753.275 -34.165 753.605 -33.835 ;
        RECT 749.195 -34.165 749.525 -33.835 ;
        RECT 747.835 -34.165 748.165 -33.835 ;
        RECT 746.475 -34.165 746.805 -33.835 ;
        RECT 745.115 -34.165 745.445 -33.835 ;
        RECT 743.755 -34.165 744.085 -33.835 ;
        RECT 742.395 -34.165 742.725 -33.835 ;
        RECT 738.315 -34.165 738.645 -33.835 ;
        RECT 734.235 -34.165 734.565 -33.835 ;
        RECT 732.875 -34.165 733.205 -33.835 ;
        RECT 731.515 -34.165 731.845 -33.835 ;
        RECT 730.155 -34.165 730.485 -33.835 ;
        RECT 728.795 -34.165 729.125 -33.835 ;
        RECT 727.435 -34.165 727.765 -33.835 ;
        RECT 721.995 -34.165 722.325 -33.835 ;
        RECT 719.275 -34.165 719.605 -33.835 ;
        RECT 717.915 -34.165 718.245 -33.835 ;
        RECT 716.555 -34.165 716.885 -33.835 ;
        RECT 715.195 -34.165 715.525 -33.835 ;
        RECT 713.835 -34.165 714.165 -33.835 ;
        RECT 712.475 -34.165 712.805 -33.835 ;
        RECT 707.035 -34.165 707.365 -33.835 ;
        RECT 704.315 -34.165 704.645 -33.835 ;
        RECT 702.955 -34.165 703.285 -33.835 ;
        RECT 701.595 -34.165 701.925 -33.835 ;
        RECT 700.235 -34.165 700.565 -33.835 ;
        RECT 698.875 -34.165 699.205 -33.835 ;
        RECT 697.515 -34.165 697.845 -33.835 ;
        RECT 692.075 -34.165 692.405 -33.835 ;
        RECT 689.355 -34.165 689.685 -33.835 ;
        RECT 687.995 -34.165 688.325 -33.835 ;
        RECT 686.635 -34.165 686.965 -33.835 ;
        RECT 685.275 -34.165 685.605 -33.835 ;
        RECT 683.915 -34.165 684.245 -33.835 ;
        RECT 682.555 -34.165 682.885 -33.835 ;
        RECT 679.835 -34.165 680.165 -33.835 ;
        RECT 677.115 -34.165 677.445 -33.835 ;
        RECT 674.395 -34.165 674.725 -33.835 ;
        RECT 673.035 -34.165 673.365 -33.835 ;
        RECT 671.675 -34.165 672.005 -33.835 ;
        RECT 670.315 -34.165 670.645 -33.835 ;
        RECT 668.955 -34.165 669.285 -33.835 ;
        RECT 667.595 -34.165 667.925 -33.835 ;
        RECT 664.875 -34.165 665.205 -33.835 ;
        RECT 662.155 -34.165 662.485 -33.835 ;
        RECT 659.435 -34.165 659.765 -33.835 ;
        RECT 658.075 -34.165 658.405 -33.835 ;
        RECT 656.715 -34.165 657.045 -33.835 ;
        RECT 655.355 -34.165 655.685 -33.835 ;
        RECT 653.995 -34.165 654.325 -33.835 ;
        RECT 652.635 -34.165 652.965 -33.835 ;
        RECT 649.915 -34.165 650.245 -33.835 ;
        RECT 647.195 -34.165 647.525 -33.835 ;
        RECT 644.475 -34.165 644.805 -33.835 ;
        RECT 643.115 -34.165 643.445 -33.835 ;
        RECT 641.755 -34.165 642.085 -33.835 ;
        RECT 640.395 -34.165 640.725 -33.835 ;
        RECT 639.035 -34.165 639.365 -33.835 ;
        RECT 637.675 -34.165 638.005 -33.835 ;
        RECT 634.955 -34.165 635.285 -33.835 ;
        RECT 632.235 -34.165 632.565 -33.835 ;
        RECT 629.515 -34.165 629.845 -33.835 ;
        RECT 628.155 -34.165 628.485 -33.835 ;
        RECT 626.795 -34.165 627.125 -33.835 ;
        RECT 625.435 -34.165 625.765 -33.835 ;
        RECT 624.075 -34.165 624.405 -33.835 ;
        RECT 622.715 -34.165 623.045 -33.835 ;
        RECT 619.995 -34.165 620.325 -33.835 ;
        RECT 617.275 -34.165 617.605 -33.835 ;
        RECT 614.555 -34.165 614.885 -33.835 ;
        RECT 613.195 -34.165 613.525 -33.835 ;
        RECT 611.835 -34.165 612.165 -33.835 ;
        RECT 610.475 -34.165 610.805 -33.835 ;
        RECT 609.115 -34.165 609.445 -33.835 ;
        RECT 607.755 -34.165 608.085 -33.835 ;
        RECT 605.035 -34.165 605.365 -33.835 ;
        RECT 602.315 -34.165 602.645 -33.835 ;
        RECT 599.595 -34.165 599.925 -33.835 ;
        RECT 598.235 -34.165 598.565 -33.835 ;
        RECT 596.875 -34.165 597.205 -33.835 ;
        RECT 595.515 -34.165 595.845 -33.835 ;
        RECT 594.155 -34.165 594.485 -33.835 ;
        RECT 592.795 -34.165 593.125 -33.835 ;
        RECT 590.075 -34.165 590.405 -33.835 ;
        RECT 587.355 -34.165 587.685 -33.835 ;
        RECT 584.635 -34.165 584.965 -33.835 ;
        RECT 583.275 -34.165 583.605 -33.835 ;
        RECT 581.915 -34.165 582.245 -33.835 ;
        RECT 580.555 -34.165 580.885 -33.835 ;
        RECT 579.195 -34.165 579.525 -33.835 ;
        RECT 577.835 -34.165 578.165 -33.835 ;
        RECT 575.115 -34.165 575.445 -33.835 ;
        RECT 572.395 -34.165 572.725 -33.835 ;
        RECT 569.675 -34.165 570.005 -33.835 ;
        RECT 568.315 -34.165 568.645 -33.835 ;
        RECT 566.955 -34.165 567.285 -33.835 ;
        RECT 565.595 -34.165 565.925 -33.835 ;
        RECT 564.235 -34.165 564.565 -33.835 ;
        RECT 562.875 -34.165 563.205 -33.835 ;
        RECT 560.155 -34.165 560.485 -33.835 ;
        RECT 557.435 -34.165 557.765 -33.835 ;
        RECT 554.715 -34.165 555.045 -33.835 ;
        RECT 553.355 -34.165 553.685 -33.835 ;
        RECT 551.995 -34.165 552.325 -33.835 ;
        RECT 550.635 -34.165 550.965 -33.835 ;
        RECT 549.275 -34.165 549.605 -33.835 ;
        RECT 547.915 -34.165 548.245 -33.835 ;
        RECT 545.195 -34.165 545.525 -33.835 ;
        RECT 542.475 -34.165 542.805 -33.835 ;
        RECT 539.755 -34.165 540.085 -33.835 ;
        RECT 538.395 -34.165 538.725 -33.835 ;
        RECT 537.035 -34.165 537.365 -33.835 ;
        RECT 535.675 -34.165 536.005 -33.835 ;
        RECT 534.315 -34.165 534.645 -33.835 ;
        RECT 532.955 -34.165 533.285 -33.835 ;
        RECT 530.235 -34.165 530.565 -33.835 ;
        RECT 527.515 -34.165 527.845 -33.835 ;
        RECT 524.795 -34.165 525.125 -33.835 ;
        RECT 523.435 -34.165 523.765 -33.835 ;
        RECT 522.075 -34.165 522.405 -33.835 ;
        RECT 520.715 -34.165 521.045 -33.835 ;
        RECT 519.355 -34.165 519.685 -33.835 ;
        RECT 517.995 -34.165 518.325 -33.835 ;
        RECT 515.275 -34.165 515.605 -33.835 ;
        RECT 512.555 -34.165 512.885 -33.835 ;
        RECT 509.835 -34.165 510.165 -33.835 ;
        RECT 508.475 -34.165 508.805 -33.835 ;
        RECT 507.115 -34.165 507.445 -33.835 ;
        RECT 505.755 -34.165 506.085 -33.835 ;
        RECT 504.395 -34.165 504.725 -33.835 ;
        RECT 500.315 -34.165 500.645 -33.835 ;
        RECT 497.595 -34.165 497.925 -33.835 ;
        RECT 494.875 -34.165 495.205 -33.835 ;
        RECT 493.515 -34.165 493.845 -33.835 ;
        RECT 492.155 -34.165 492.485 -33.835 ;
        RECT 490.795 -34.165 491.125 -33.835 ;
        RECT 489.435 -34.165 489.765 -33.835 ;
        RECT 485.355 -34.165 485.685 -33.835 ;
        RECT 482.635 -34.165 482.965 -33.835 ;
        RECT 479.915 -34.165 480.245 -33.835 ;
        RECT 478.555 -34.165 478.885 -33.835 ;
        RECT 477.195 -34.165 477.525 -33.835 ;
        RECT 475.835 -34.165 476.165 -33.835 ;
        RECT 474.475 -34.165 474.805 -33.835 ;
        RECT 470.395 -34.165 470.725 -33.835 ;
        RECT 467.675 -34.165 468.005 -33.835 ;
        RECT 464.955 -34.165 465.285 -33.835 ;
        RECT 463.595 -34.165 463.925 -33.835 ;
        RECT 462.235 -34.165 462.565 -33.835 ;
        RECT 460.875 -34.165 461.205 -33.835 ;
        RECT 459.515 -34.165 459.845 -33.835 ;
        RECT 455.435 -34.165 455.765 -33.835 ;
        RECT 452.715 -34.165 453.045 -33.835 ;
        RECT 449.995 -34.165 450.325 -33.835 ;
        RECT 448.635 -34.165 448.965 -33.835 ;
        RECT 447.275 -34.165 447.605 -33.835 ;
        RECT 445.915 -34.165 446.245 -33.835 ;
        RECT 444.555 -34.165 444.885 -33.835 ;
        RECT 440.475 -34.165 440.805 -33.835 ;
        RECT 436.395 -34.165 436.725 -33.835 ;
        RECT 435.035 -34.165 435.365 -33.835 ;
        RECT 433.675 -34.165 434.005 -33.835 ;
        RECT 432.315 -34.165 432.645 -33.835 ;
        RECT 430.955 -34.165 431.285 -33.835 ;
        RECT 429.595 -34.165 429.925 -33.835 ;
        RECT 425.515 -34.165 425.845 -33.835 ;
        RECT 421.435 -34.165 421.765 -33.835 ;
        RECT 420.075 -34.165 420.405 -33.835 ;
        RECT 418.715 -34.165 419.045 -33.835 ;
        RECT 417.355 -34.165 417.685 -33.835 ;
        RECT 415.995 -34.165 416.325 -33.835 ;
        RECT 414.635 -34.165 414.965 -33.835 ;
        RECT 410.555 -34.165 410.885 -33.835 ;
        RECT 406.475 -34.165 406.805 -33.835 ;
        RECT 405.115 -34.165 405.445 -33.835 ;
        RECT 403.755 -34.165 404.085 -33.835 ;
        RECT 402.395 -34.165 402.725 -33.835 ;
        RECT 401.035 -34.165 401.365 -33.835 ;
        RECT 399.675 -34.165 400.005 -33.835 ;
        RECT 395.595 -34.165 395.925 -33.835 ;
        RECT 394.235 -34.165 394.565 -33.835 ;
        RECT 391.515 -34.165 391.845 -33.835 ;
        RECT 390.155 -34.165 390.485 -33.835 ;
        RECT 388.795 -34.165 389.125 -33.835 ;
        RECT 387.435 -34.165 387.765 -33.835 ;
        RECT 386.075 -34.165 386.405 -33.835 ;
        RECT 384.715 -34.165 385.045 -33.835 ;
        RECT 379.275 -34.165 379.605 -33.835 ;
        RECT 376.555 -34.165 376.885 -33.835 ;
        RECT 375.195 -34.165 375.525 -33.835 ;
        RECT 373.835 -34.165 374.165 -33.835 ;
        RECT 372.475 -34.165 372.805 -33.835 ;
        RECT 371.115 -34.165 371.445 -33.835 ;
        RECT 369.755 -34.165 370.085 -33.835 ;
        RECT 364.315 -34.165 364.645 -33.835 ;
        RECT 361.595 -34.165 361.925 -33.835 ;
        RECT 360.235 -34.165 360.565 -33.835 ;
        RECT 358.875 -34.165 359.205 -33.835 ;
        RECT 357.515 -34.165 357.845 -33.835 ;
        RECT 356.155 -34.165 356.485 -33.835 ;
        RECT 354.795 -34.165 355.125 -33.835 ;
        RECT 349.355 -34.165 349.685 -33.835 ;
        RECT 346.635 -34.165 346.965 -33.835 ;
        RECT 345.275 -34.165 345.605 -33.835 ;
        RECT 343.915 -34.165 344.245 -33.835 ;
        RECT 342.555 -34.165 342.885 -33.835 ;
        RECT 341.195 -34.165 341.525 -33.835 ;
        RECT 339.835 -34.165 340.165 -33.835 ;
        RECT 337.115 -34.165 337.445 -33.835 ;
        RECT 334.395 -34.165 334.725 -33.835 ;
        RECT 331.675 -34.165 332.005 -33.835 ;
        RECT 330.315 -34.165 330.645 -33.835 ;
        RECT 328.955 -34.165 329.285 -33.835 ;
        RECT 327.595 -34.165 327.925 -33.835 ;
        RECT 326.235 -34.165 326.565 -33.835 ;
        RECT 324.875 -34.165 325.205 -33.835 ;
        RECT 322.155 -34.165 322.485 -33.835 ;
        RECT 319.435 -34.165 319.765 -33.835 ;
        RECT 316.715 -34.165 317.045 -33.835 ;
        RECT 315.355 -34.165 315.685 -33.835 ;
        RECT 313.995 -34.165 314.325 -33.835 ;
        RECT 312.635 -34.165 312.965 -33.835 ;
        RECT 311.275 -34.165 311.605 -33.835 ;
        RECT 309.915 -34.165 310.245 -33.835 ;
        RECT 307.195 -34.165 307.525 -33.835 ;
        RECT 304.475 -34.165 304.805 -33.835 ;
        RECT 301.755 -34.165 302.085 -33.835 ;
        RECT 300.395 -34.165 300.725 -33.835 ;
        RECT 299.035 -34.165 299.365 -33.835 ;
        RECT 297.675 -34.165 298.005 -33.835 ;
        RECT 296.315 -34.165 296.645 -33.835 ;
        RECT 294.955 -34.165 295.285 -33.835 ;
        RECT 292.235 -34.165 292.565 -33.835 ;
        RECT 289.515 -34.165 289.845 -33.835 ;
        RECT 286.795 -34.165 287.125 -33.835 ;
        RECT 285.435 -34.165 285.765 -33.835 ;
        RECT 284.075 -34.165 284.405 -33.835 ;
        RECT 282.715 -34.165 283.045 -33.835 ;
        RECT 281.355 -34.165 281.685 -33.835 ;
        RECT 279.995 -34.165 280.325 -33.835 ;
        RECT 277.275 -34.165 277.605 -33.835 ;
        RECT 274.555 -34.165 274.885 -33.835 ;
        RECT 271.835 -34.165 272.165 -33.835 ;
        RECT 270.475 -34.165 270.805 -33.835 ;
        RECT 269.115 -34.165 269.445 -33.835 ;
        RECT 267.755 -34.165 268.085 -33.835 ;
        RECT 266.395 -34.165 266.725 -33.835 ;
        RECT 265.035 -34.165 265.365 -33.835 ;
        RECT 262.315 -34.165 262.645 -33.835 ;
        RECT 259.595 -34.165 259.925 -33.835 ;
        RECT 256.875 -34.165 257.205 -33.835 ;
        RECT 255.515 -34.165 255.845 -33.835 ;
        RECT 254.155 -34.165 254.485 -33.835 ;
        RECT 252.795 -34.165 253.125 -33.835 ;
        RECT 251.435 -34.165 251.765 -33.835 ;
        RECT 250.075 -34.165 250.405 -33.835 ;
        RECT 247.355 -34.165 247.685 -33.835 ;
        RECT 244.635 -34.165 244.965 -33.835 ;
        RECT 241.915 -34.165 242.245 -33.835 ;
        RECT 240.555 -34.165 240.885 -33.835 ;
        RECT 239.195 -34.165 239.525 -33.835 ;
        RECT 237.835 -34.165 238.165 -33.835 ;
        RECT 236.475 -34.165 236.805 -33.835 ;
        RECT 235.115 -34.165 235.445 -33.835 ;
        RECT 232.395 -34.165 232.725 -33.835 ;
        RECT 229.675 -34.165 230.005 -33.835 ;
        RECT 226.955 -34.165 227.285 -33.835 ;
        RECT 225.595 -34.165 225.925 -33.835 ;
        RECT 224.235 -34.165 224.565 -33.835 ;
        RECT 222.875 -34.165 223.205 -33.835 ;
        RECT 221.515 -34.165 221.845 -33.835 ;
        RECT 220.155 -34.165 220.485 -33.835 ;
        RECT 217.435 -34.165 217.765 -33.835 ;
        RECT 214.715 -34.165 215.045 -33.835 ;
        RECT 211.995 -34.165 212.325 -33.835 ;
        RECT 210.635 -34.165 210.965 -33.835 ;
        RECT 209.275 -34.165 209.605 -33.835 ;
        RECT 207.915 -34.165 208.245 -33.835 ;
        RECT 206.555 -34.165 206.885 -33.835 ;
        RECT 205.195 -34.165 205.525 -33.835 ;
        RECT 202.475 -34.165 202.805 -33.835 ;
        RECT 199.755 -34.165 200.085 -33.835 ;
        RECT 197.035 -34.165 197.365 -33.835 ;
        RECT 195.675 -34.165 196.005 -33.835 ;
        RECT 194.315 -34.165 194.645 -33.835 ;
        RECT 192.955 -34.165 193.285 -33.835 ;
        RECT 191.595 -34.165 191.925 -33.835 ;
        RECT 190.235 -34.165 190.565 -33.835 ;
        RECT 187.515 -34.165 187.845 -33.835 ;
        RECT 184.795 -34.165 185.125 -33.835 ;
        RECT 182.075 -34.165 182.405 -33.835 ;
        RECT 180.715 -34.165 181.045 -33.835 ;
        RECT 179.355 -34.165 179.685 -33.835 ;
        RECT 177.995 -34.165 178.325 -33.835 ;
        RECT 176.635 -34.165 176.965 -33.835 ;
        RECT 175.275 -34.165 175.605 -33.835 ;
        RECT 172.555 -34.165 172.885 -33.835 ;
        RECT 169.835 -34.165 170.165 -33.835 ;
        RECT 167.115 -34.165 167.445 -33.835 ;
        RECT 165.755 -34.165 166.085 -33.835 ;
        RECT 164.395 -34.165 164.725 -33.835 ;
        RECT 163.035 -34.165 163.365 -33.835 ;
        RECT 161.675 -34.165 162.005 -33.835 ;
        RECT 157.595 -34.165 157.925 -33.835 ;
        RECT 154.875 -34.165 155.205 -33.835 ;
        RECT 152.155 -34.165 152.485 -33.835 ;
        RECT 150.795 -34.165 151.125 -33.835 ;
        RECT 149.435 -34.165 149.765 -33.835 ;
        RECT 148.075 -34.165 148.405 -33.835 ;
        RECT 146.715 -34.165 147.045 -33.835 ;
        RECT 142.635 -34.165 142.965 -33.835 ;
        RECT 139.915 -34.165 140.245 -33.835 ;
        RECT 137.195 -34.165 137.525 -33.835 ;
        RECT 135.835 -34.165 136.165 -33.835 ;
        RECT 134.475 -34.165 134.805 -33.835 ;
        RECT 133.115 -34.165 133.445 -33.835 ;
        RECT 131.755 -34.165 132.085 -33.835 ;
        RECT 127.675 -34.165 128.005 -33.835 ;
        RECT 124.955 -34.165 125.285 -33.835 ;
        RECT 122.235 -34.165 122.565 -33.835 ;
        RECT 120.875 -34.165 121.205 -33.835 ;
        RECT 119.515 -34.165 119.845 -33.835 ;
        RECT 118.155 -34.165 118.485 -33.835 ;
        RECT 116.795 -34.165 117.125 -33.835 ;
        RECT 112.715 -34.165 113.045 -33.835 ;
        RECT 109.995 -34.165 110.325 -33.835 ;
        RECT 107.275 -34.165 107.605 -33.835 ;
        RECT 105.915 -34.165 106.245 -33.835 ;
        RECT 104.555 -34.165 104.885 -33.835 ;
        RECT 103.195 -34.165 103.525 -33.835 ;
        RECT 101.835 -34.165 102.165 -33.835 ;
        RECT 97.755 -34.165 98.085 -33.835 ;
        RECT 93.675 -34.165 94.005 -33.835 ;
        RECT 92.315 -34.165 92.645 -33.835 ;
        RECT 90.955 -34.165 91.285 -33.835 ;
        RECT 89.595 -34.165 89.925 -33.835 ;
        RECT 88.235 -34.165 88.565 -33.835 ;
        RECT 86.875 -34.165 87.205 -33.835 ;
        RECT 82.795 -34.165 83.125 -33.835 ;
        RECT 78.715 -34.165 79.045 -33.835 ;
        RECT 77.355 -34.165 77.685 -33.835 ;
        RECT 75.995 -34.165 76.325 -33.835 ;
        RECT 74.635 -34.165 74.965 -33.835 ;
        RECT 73.275 -34.165 73.605 -33.835 ;
        RECT 71.915 -34.165 72.245 -33.835 ;
        RECT 67.835 -34.165 68.165 -33.835 ;
        RECT 63.755 -34.165 64.085 -33.835 ;
        RECT 62.395 -34.165 62.725 -33.835 ;
        RECT 61.035 -34.165 61.365 -33.835 ;
        RECT 59.675 -34.165 60.005 -33.835 ;
        RECT 58.315 -34.165 58.645 -33.835 ;
        RECT 56.955 -34.165 57.285 -33.835 ;
        RECT 51.515 -34.165 51.845 -33.835 ;
        RECT 48.795 -34.165 49.125 -33.835 ;
        RECT 47.435 -34.165 47.765 -33.835 ;
        RECT 46.075 -34.165 46.405 -33.835 ;
        RECT 44.715 -34.165 45.045 -33.835 ;
        RECT 43.355 -34.165 43.685 -33.835 ;
        RECT 41.995 -34.165 42.325 -33.835 ;
        RECT 36.555 -34.165 36.885 -33.835 ;
        RECT 33.835 -34.165 34.165 -33.835 ;
        RECT 32.475 -34.165 32.805 -33.835 ;
        RECT 31.115 -34.165 31.445 -33.835 ;
        RECT 29.755 -34.165 30.085 -33.835 ;
        RECT 28.395 -34.165 28.725 -33.835 ;
        RECT 27.035 -34.165 27.365 -33.835 ;
        RECT 21.595 -34.165 21.925 -33.835 ;
        RECT 18.875 -34.165 19.205 -33.835 ;
        RECT 17.515 -34.165 17.845 -33.835 ;
        RECT 16.155 -34.165 16.485 -33.835 ;
        RECT 14.795 -34.165 15.125 -33.835 ;
        RECT 13.435 -34.165 13.765 -33.835 ;
        RECT 12.075 -34.165 12.405 -33.835 ;
        RECT 10.715 -34.165 11.045 -33.835 ;
        RECT 7.995 -34.165 8.325 -33.835 ;
        RECT 6.635 -34.165 6.965 -33.835 ;
        RECT 5.275 -34.165 5.605 -33.835 ;
        RECT 3.915 -34.165 4.245 -33.835 ;
        RECT 2.555 -34.165 2.885 -33.835 ;
        RECT 1.195 -34.165 1.525 -33.835 ;
        RECT -0.165 -34.165 0.165 -33.835 ;
        RECT -1.525 -34.165 -1.195 -33.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -35.525 954.885 -35.195 ;
        RECT 949.12 -35.52 954.885 -35.2 ;
        RECT 953.195 -35.525 953.525 -35.195 ;
        RECT 951.835 -35.525 952.165 -35.195 ;
        RECT 950.475 -35.525 950.805 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -23.285 954.885 -22.955 ;
        RECT 945.035 -23.28 954.885 -22.96 ;
        RECT 953.195 -23.285 953.525 -22.955 ;
        RECT 951.835 -23.285 952.165 -22.955 ;
        RECT 950.475 -23.285 950.805 -22.955 ;
        RECT 946.395 -23.285 946.725 -22.955 ;
        RECT 945.035 -23.285 945.365 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -26.005 954.885 -25.675 ;
        RECT 934.84 -26 954.885 -25.68 ;
        RECT 953.195 -26.005 953.525 -25.675 ;
        RECT 951.835 -26.005 952.165 -25.675 ;
        RECT 950.475 -26.005 950.805 -25.675 ;
        RECT 946.395 -26.005 946.725 -25.675 ;
        RECT 945.035 -26.005 945.365 -25.675 ;
        RECT 943.675 -26.005 944.005 -25.675 ;
        RECT 942.315 -26.005 942.645 -25.675 ;
        RECT 940.955 -26.005 941.285 -25.675 ;
        RECT 939.595 -26.005 939.925 -25.675 ;
        RECT 938.235 -26.005 938.565 -25.675 ;
        RECT 936.875 -26.005 937.205 -25.675 ;
        RECT 935.515 -26.005 935.845 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -27.365 954.885 -27.035 ;
        RECT 930.76 -27.36 954.885 -27.04 ;
        RECT 953.195 -27.365 953.525 -27.035 ;
        RECT 951.835 -27.365 952.165 -27.035 ;
        RECT 950.475 -27.365 950.805 -27.035 ;
        RECT 946.395 -27.365 946.725 -27.035 ;
        RECT 945.035 -27.365 945.365 -27.035 ;
        RECT 943.675 -27.365 944.005 -27.035 ;
        RECT 942.315 -27.365 942.645 -27.035 ;
        RECT 940.955 -27.365 941.285 -27.035 ;
        RECT 939.595 -27.365 939.925 -27.035 ;
        RECT 938.235 -27.365 938.565 -27.035 ;
        RECT 936.875 -27.365 937.205 -27.035 ;
        RECT 935.515 -27.365 935.845 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -28.725 954.885 -28.395 ;
        RECT -1.525 -28.72 954.885 -28.4 ;
        RECT 953.195 -28.725 953.525 -28.395 ;
        RECT 951.835 -28.725 952.165 -28.395 ;
        RECT 950.475 -28.725 950.805 -28.395 ;
        RECT 946.395 -28.725 946.725 -28.395 ;
        RECT 945.035 -28.725 945.365 -28.395 ;
        RECT 943.675 -28.725 944.005 -28.395 ;
        RECT 942.315 -28.725 942.645 -28.395 ;
        RECT 940.955 -28.725 941.285 -28.395 ;
        RECT 939.595 -28.725 939.925 -28.395 ;
        RECT 938.235 -28.725 938.565 -28.395 ;
        RECT 936.875 -28.725 937.205 -28.395 ;
        RECT 935.515 -28.725 935.845 -28.395 ;
        RECT 930.075 -28.725 930.405 -28.395 ;
        RECT 928.715 -28.725 929.045 -28.395 ;
        RECT 924.635 -28.725 924.965 -28.395 ;
        RECT 923.275 -28.725 923.605 -28.395 ;
        RECT 921.915 -28.725 922.245 -28.395 ;
        RECT 920.555 -28.725 920.885 -28.395 ;
        RECT 915.115 -28.725 915.445 -28.395 ;
        RECT 913.755 -28.725 914.085 -28.395 ;
        RECT 909.675 -28.725 910.005 -28.395 ;
        RECT 908.315 -28.725 908.645 -28.395 ;
        RECT 906.955 -28.725 907.285 -28.395 ;
        RECT 905.595 -28.725 905.925 -28.395 ;
        RECT 900.155 -28.725 900.485 -28.395 ;
        RECT 898.795 -28.725 899.125 -28.395 ;
        RECT 894.715 -28.725 895.045 -28.395 ;
        RECT 893.355 -28.725 893.685 -28.395 ;
        RECT 891.995 -28.725 892.325 -28.395 ;
        RECT 890.635 -28.725 890.965 -28.395 ;
        RECT 885.195 -28.725 885.525 -28.395 ;
        RECT 883.835 -28.725 884.165 -28.395 ;
        RECT 879.755 -28.725 880.085 -28.395 ;
        RECT 878.395 -28.725 878.725 -28.395 ;
        RECT 877.035 -28.725 877.365 -28.395 ;
        RECT 875.675 -28.725 876.005 -28.395 ;
        RECT 870.235 -28.725 870.565 -28.395 ;
        RECT 868.875 -28.725 869.205 -28.395 ;
        RECT 864.795 -28.725 865.125 -28.395 ;
        RECT 863.435 -28.725 863.765 -28.395 ;
        RECT 862.075 -28.725 862.405 -28.395 ;
        RECT 860.715 -28.725 861.045 -28.395 ;
        RECT 857.995 -28.725 858.325 -28.395 ;
        RECT 855.275 -28.725 855.605 -28.395 ;
        RECT 853.915 -28.725 854.245 -28.395 ;
        RECT 849.835 -28.725 850.165 -28.395 ;
        RECT 848.475 -28.725 848.805 -28.395 ;
        RECT 847.115 -28.725 847.445 -28.395 ;
        RECT 845.755 -28.725 846.085 -28.395 ;
        RECT 843.035 -28.725 843.365 -28.395 ;
        RECT 840.315 -28.725 840.645 -28.395 ;
        RECT 838.955 -28.725 839.285 -28.395 ;
        RECT 834.875 -28.725 835.205 -28.395 ;
        RECT 833.515 -28.725 833.845 -28.395 ;
        RECT 832.155 -28.725 832.485 -28.395 ;
        RECT 828.075 -28.725 828.405 -28.395 ;
        RECT 825.355 -28.725 825.685 -28.395 ;
        RECT 823.995 -28.725 824.325 -28.395 ;
        RECT 819.915 -28.725 820.245 -28.395 ;
        RECT 818.555 -28.725 818.885 -28.395 ;
        RECT 817.195 -28.725 817.525 -28.395 ;
        RECT 813.115 -28.725 813.445 -28.395 ;
        RECT 810.395 -28.725 810.725 -28.395 ;
        RECT 804.955 -28.725 805.285 -28.395 ;
        RECT 803.595 -28.725 803.925 -28.395 ;
        RECT 802.235 -28.725 802.565 -28.395 ;
        RECT 798.155 -28.725 798.485 -28.395 ;
        RECT 795.435 -28.725 795.765 -28.395 ;
        RECT 791.355 -28.725 791.685 -28.395 ;
        RECT 789.995 -28.725 790.325 -28.395 ;
        RECT 788.635 -28.725 788.965 -28.395 ;
        RECT 787.275 -28.725 787.605 -28.395 ;
        RECT 783.195 -28.725 783.525 -28.395 ;
        RECT 780.475 -28.725 780.805 -28.395 ;
        RECT 776.395 -28.725 776.725 -28.395 ;
        RECT 775.035 -28.725 775.365 -28.395 ;
        RECT 773.675 -28.725 774.005 -28.395 ;
        RECT 772.315 -28.725 772.645 -28.395 ;
        RECT 768.235 -28.725 768.565 -28.395 ;
        RECT 761.435 -28.725 761.765 -28.395 ;
        RECT 760.075 -28.725 760.405 -28.395 ;
        RECT 758.715 -28.725 759.045 -28.395 ;
        RECT 757.355 -28.725 757.685 -28.395 ;
        RECT 753.275 -28.725 753.605 -28.395 ;
        RECT 750.555 -28.725 750.885 -28.395 ;
        RECT 746.475 -28.725 746.805 -28.395 ;
        RECT 745.115 -28.725 745.445 -28.395 ;
        RECT 743.755 -28.725 744.085 -28.395 ;
        RECT 742.395 -28.725 742.725 -28.395 ;
        RECT 738.315 -28.725 738.645 -28.395 ;
        RECT 735.595 -28.725 735.925 -28.395 ;
        RECT 731.515 -28.725 731.845 -28.395 ;
        RECT 730.155 -28.725 730.485 -28.395 ;
        RECT 728.795 -28.725 729.125 -28.395 ;
        RECT 727.435 -28.725 727.765 -28.395 ;
        RECT 721.995 -28.725 722.325 -28.395 ;
        RECT 720.635 -28.725 720.965 -28.395 ;
        RECT 716.555 -28.725 716.885 -28.395 ;
        RECT 715.195 -28.725 715.525 -28.395 ;
        RECT 713.835 -28.725 714.165 -28.395 ;
        RECT 712.475 -28.725 712.805 -28.395 ;
        RECT 707.035 -28.725 707.365 -28.395 ;
        RECT 705.675 -28.725 706.005 -28.395 ;
        RECT 701.595 -28.725 701.925 -28.395 ;
        RECT 700.235 -28.725 700.565 -28.395 ;
        RECT 698.875 -28.725 699.205 -28.395 ;
        RECT 697.515 -28.725 697.845 -28.395 ;
        RECT 692.075 -28.725 692.405 -28.395 ;
        RECT 690.715 -28.725 691.045 -28.395 ;
        RECT 686.635 -28.725 686.965 -28.395 ;
        RECT 685.275 -28.725 685.605 -28.395 ;
        RECT 683.915 -28.725 684.245 -28.395 ;
        RECT 682.555 -28.725 682.885 -28.395 ;
        RECT 677.115 -28.725 677.445 -28.395 ;
        RECT 675.755 -28.725 676.085 -28.395 ;
        RECT 671.675 -28.725 672.005 -28.395 ;
        RECT 670.315 -28.725 670.645 -28.395 ;
        RECT 668.955 -28.725 669.285 -28.395 ;
        RECT 667.595 -28.725 667.925 -28.395 ;
        RECT 662.155 -28.725 662.485 -28.395 ;
        RECT 660.795 -28.725 661.125 -28.395 ;
        RECT 656.715 -28.725 657.045 -28.395 ;
        RECT 655.355 -28.725 655.685 -28.395 ;
        RECT 653.995 -28.725 654.325 -28.395 ;
        RECT 652.635 -28.725 652.965 -28.395 ;
        RECT 647.195 -28.725 647.525 -28.395 ;
        RECT 645.835 -28.725 646.165 -28.395 ;
        RECT 641.755 -28.725 642.085 -28.395 ;
        RECT 640.395 -28.725 640.725 -28.395 ;
        RECT 639.035 -28.725 639.365 -28.395 ;
        RECT 637.675 -28.725 638.005 -28.395 ;
        RECT 632.235 -28.725 632.565 -28.395 ;
        RECT 630.875 -28.725 631.205 -28.395 ;
        RECT 626.795 -28.725 627.125 -28.395 ;
        RECT 625.435 -28.725 625.765 -28.395 ;
        RECT 624.075 -28.725 624.405 -28.395 ;
        RECT 622.715 -28.725 623.045 -28.395 ;
        RECT 617.275 -28.725 617.605 -28.395 ;
        RECT 615.915 -28.725 616.245 -28.395 ;
        RECT 611.835 -28.725 612.165 -28.395 ;
        RECT 610.475 -28.725 610.805 -28.395 ;
        RECT 609.115 -28.725 609.445 -28.395 ;
        RECT 607.755 -28.725 608.085 -28.395 ;
        RECT 602.315 -28.725 602.645 -28.395 ;
        RECT 600.955 -28.725 601.285 -28.395 ;
        RECT 596.875 -28.725 597.205 -28.395 ;
        RECT 595.515 -28.725 595.845 -28.395 ;
        RECT 594.155 -28.725 594.485 -28.395 ;
        RECT 592.795 -28.725 593.125 -28.395 ;
        RECT 587.355 -28.725 587.685 -28.395 ;
        RECT 585.995 -28.725 586.325 -28.395 ;
        RECT 581.915 -28.725 582.245 -28.395 ;
        RECT 580.555 -28.725 580.885 -28.395 ;
        RECT 579.195 -28.725 579.525 -28.395 ;
        RECT 577.835 -28.725 578.165 -28.395 ;
        RECT 572.395 -28.725 572.725 -28.395 ;
        RECT 571.035 -28.725 571.365 -28.395 ;
        RECT 566.955 -28.725 567.285 -28.395 ;
        RECT 565.595 -28.725 565.925 -28.395 ;
        RECT 564.235 -28.725 564.565 -28.395 ;
        RECT 562.875 -28.725 563.205 -28.395 ;
        RECT 557.435 -28.725 557.765 -28.395 ;
        RECT 556.075 -28.725 556.405 -28.395 ;
        RECT 551.995 -28.725 552.325 -28.395 ;
        RECT 550.635 -28.725 550.965 -28.395 ;
        RECT 549.275 -28.725 549.605 -28.395 ;
        RECT 547.915 -28.725 548.245 -28.395 ;
        RECT 542.475 -28.725 542.805 -28.395 ;
        RECT 541.115 -28.725 541.445 -28.395 ;
        RECT 537.035 -28.725 537.365 -28.395 ;
        RECT 535.675 -28.725 536.005 -28.395 ;
        RECT 534.315 -28.725 534.645 -28.395 ;
        RECT 532.955 -28.725 533.285 -28.395 ;
        RECT 527.515 -28.725 527.845 -28.395 ;
        RECT 526.155 -28.725 526.485 -28.395 ;
        RECT 522.075 -28.725 522.405 -28.395 ;
        RECT 520.715 -28.725 521.045 -28.395 ;
        RECT 519.355 -28.725 519.685 -28.395 ;
        RECT 517.995 -28.725 518.325 -28.395 ;
        RECT 515.275 -28.725 515.605 -28.395 ;
        RECT 512.555 -28.725 512.885 -28.395 ;
        RECT 511.195 -28.725 511.525 -28.395 ;
        RECT 507.115 -28.725 507.445 -28.395 ;
        RECT 505.755 -28.725 506.085 -28.395 ;
        RECT 504.395 -28.725 504.725 -28.395 ;
        RECT 500.315 -28.725 500.645 -28.395 ;
        RECT 497.595 -28.725 497.925 -28.395 ;
        RECT 496.235 -28.725 496.565 -28.395 ;
        RECT 492.155 -28.725 492.485 -28.395 ;
        RECT 490.795 -28.725 491.125 -28.395 ;
        RECT 489.435 -28.725 489.765 -28.395 ;
        RECT 485.355 -28.725 485.685 -28.395 ;
        RECT 482.635 -28.725 482.965 -28.395 ;
        RECT 481.275 -28.725 481.605 -28.395 ;
        RECT 477.195 -28.725 477.525 -28.395 ;
        RECT 475.835 -28.725 476.165 -28.395 ;
        RECT 474.475 -28.725 474.805 -28.395 ;
        RECT 470.395 -28.725 470.725 -28.395 ;
        RECT 467.675 -28.725 468.005 -28.395 ;
        RECT 463.595 -28.725 463.925 -28.395 ;
        RECT 462.235 -28.725 462.565 -28.395 ;
        RECT 460.875 -28.725 461.205 -28.395 ;
        RECT 459.515 -28.725 459.845 -28.395 ;
        RECT 455.435 -28.725 455.765 -28.395 ;
        RECT 452.715 -28.725 453.045 -28.395 ;
        RECT 448.635 -28.725 448.965 -28.395 ;
        RECT 447.275 -28.725 447.605 -28.395 ;
        RECT 445.915 -28.725 446.245 -28.395 ;
        RECT 444.555 -28.725 444.885 -28.395 ;
        RECT 440.475 -28.725 440.805 -28.395 ;
        RECT 433.675 -28.725 434.005 -28.395 ;
        RECT 432.315 -28.725 432.645 -28.395 ;
        RECT 430.955 -28.725 431.285 -28.395 ;
        RECT 429.595 -28.725 429.925 -28.395 ;
        RECT 425.515 -28.725 425.845 -28.395 ;
        RECT 418.715 -28.725 419.045 -28.395 ;
        RECT 417.355 -28.725 417.685 -28.395 ;
        RECT 415.995 -28.725 416.325 -28.395 ;
        RECT 414.635 -28.725 414.965 -28.395 ;
        RECT 410.555 -28.725 410.885 -28.395 ;
        RECT 407.835 -28.725 408.165 -28.395 ;
        RECT 403.755 -28.725 404.085 -28.395 ;
        RECT 402.395 -28.725 402.725 -28.395 ;
        RECT 401.035 -28.725 401.365 -28.395 ;
        RECT 399.675 -28.725 400.005 -28.395 ;
        RECT 395.595 -28.725 395.925 -28.395 ;
        RECT 394.235 -28.725 394.565 -28.395 ;
        RECT 392.875 -28.725 393.205 -28.395 ;
        RECT 388.795 -28.725 389.125 -28.395 ;
        RECT 387.435 -28.725 387.765 -28.395 ;
        RECT 386.075 -28.725 386.405 -28.395 ;
        RECT 384.715 -28.725 385.045 -28.395 ;
        RECT 379.275 -28.725 379.605 -28.395 ;
        RECT 377.915 -28.725 378.245 -28.395 ;
        RECT 373.835 -28.725 374.165 -28.395 ;
        RECT 372.475 -28.725 372.805 -28.395 ;
        RECT 371.115 -28.725 371.445 -28.395 ;
        RECT 369.755 -28.725 370.085 -28.395 ;
        RECT 364.315 -28.725 364.645 -28.395 ;
        RECT 362.955 -28.725 363.285 -28.395 ;
        RECT 358.875 -28.725 359.205 -28.395 ;
        RECT 357.515 -28.725 357.845 -28.395 ;
        RECT 356.155 -28.725 356.485 -28.395 ;
        RECT 354.795 -28.725 355.125 -28.395 ;
        RECT 349.355 -28.725 349.685 -28.395 ;
        RECT 347.995 -28.725 348.325 -28.395 ;
        RECT 343.915 -28.725 344.245 -28.395 ;
        RECT 342.555 -28.725 342.885 -28.395 ;
        RECT 341.195 -28.725 341.525 -28.395 ;
        RECT 339.835 -28.725 340.165 -28.395 ;
        RECT 334.395 -28.725 334.725 -28.395 ;
        RECT 333.035 -28.725 333.365 -28.395 ;
        RECT 328.955 -28.725 329.285 -28.395 ;
        RECT 327.595 -28.725 327.925 -28.395 ;
        RECT 326.235 -28.725 326.565 -28.395 ;
        RECT 324.875 -28.725 325.205 -28.395 ;
        RECT 319.435 -28.725 319.765 -28.395 ;
        RECT 318.075 -28.725 318.405 -28.395 ;
        RECT 313.995 -28.725 314.325 -28.395 ;
        RECT 312.635 -28.725 312.965 -28.395 ;
        RECT 311.275 -28.725 311.605 -28.395 ;
        RECT 309.915 -28.725 310.245 -28.395 ;
        RECT 304.475 -28.725 304.805 -28.395 ;
        RECT 303.115 -28.725 303.445 -28.395 ;
        RECT 299.035 -28.725 299.365 -28.395 ;
        RECT 297.675 -28.725 298.005 -28.395 ;
        RECT 296.315 -28.725 296.645 -28.395 ;
        RECT 294.955 -28.725 295.285 -28.395 ;
        RECT 289.515 -28.725 289.845 -28.395 ;
        RECT 288.155 -28.725 288.485 -28.395 ;
        RECT 284.075 -28.725 284.405 -28.395 ;
        RECT 282.715 -28.725 283.045 -28.395 ;
        RECT 281.355 -28.725 281.685 -28.395 ;
        RECT 279.995 -28.725 280.325 -28.395 ;
        RECT 274.555 -28.725 274.885 -28.395 ;
        RECT 273.195 -28.725 273.525 -28.395 ;
        RECT 269.115 -28.725 269.445 -28.395 ;
        RECT 267.755 -28.725 268.085 -28.395 ;
        RECT 266.395 -28.725 266.725 -28.395 ;
        RECT 265.035 -28.725 265.365 -28.395 ;
        RECT 259.595 -28.725 259.925 -28.395 ;
        RECT 258.235 -28.725 258.565 -28.395 ;
        RECT 254.155 -28.725 254.485 -28.395 ;
        RECT 252.795 -28.725 253.125 -28.395 ;
        RECT 251.435 -28.725 251.765 -28.395 ;
        RECT 250.075 -28.725 250.405 -28.395 ;
        RECT 244.635 -28.725 244.965 -28.395 ;
        RECT 243.275 -28.725 243.605 -28.395 ;
        RECT 239.195 -28.725 239.525 -28.395 ;
        RECT 237.835 -28.725 238.165 -28.395 ;
        RECT 236.475 -28.725 236.805 -28.395 ;
        RECT 235.115 -28.725 235.445 -28.395 ;
        RECT 229.675 -28.725 230.005 -28.395 ;
        RECT 228.315 -28.725 228.645 -28.395 ;
        RECT 224.235 -28.725 224.565 -28.395 ;
        RECT 222.875 -28.725 223.205 -28.395 ;
        RECT 221.515 -28.725 221.845 -28.395 ;
        RECT 220.155 -28.725 220.485 -28.395 ;
        RECT 214.715 -28.725 215.045 -28.395 ;
        RECT 213.355 -28.725 213.685 -28.395 ;
        RECT 209.275 -28.725 209.605 -28.395 ;
        RECT 207.915 -28.725 208.245 -28.395 ;
        RECT 206.555 -28.725 206.885 -28.395 ;
        RECT 205.195 -28.725 205.525 -28.395 ;
        RECT 199.755 -28.725 200.085 -28.395 ;
        RECT 198.395 -28.725 198.725 -28.395 ;
        RECT 194.315 -28.725 194.645 -28.395 ;
        RECT 192.955 -28.725 193.285 -28.395 ;
        RECT 191.595 -28.725 191.925 -28.395 ;
        RECT 190.235 -28.725 190.565 -28.395 ;
        RECT 184.795 -28.725 185.125 -28.395 ;
        RECT 183.435 -28.725 183.765 -28.395 ;
        RECT 179.355 -28.725 179.685 -28.395 ;
        RECT 177.995 -28.725 178.325 -28.395 ;
        RECT 176.635 -28.725 176.965 -28.395 ;
        RECT 175.275 -28.725 175.605 -28.395 ;
        RECT 172.555 -28.725 172.885 -28.395 ;
        RECT 169.835 -28.725 170.165 -28.395 ;
        RECT 168.475 -28.725 168.805 -28.395 ;
        RECT 164.395 -28.725 164.725 -28.395 ;
        RECT 163.035 -28.725 163.365 -28.395 ;
        RECT 161.675 -28.725 162.005 -28.395 ;
        RECT 157.595 -28.725 157.925 -28.395 ;
        RECT 154.875 -28.725 155.205 -28.395 ;
        RECT 153.515 -28.725 153.845 -28.395 ;
        RECT 149.435 -28.725 149.765 -28.395 ;
        RECT 148.075 -28.725 148.405 -28.395 ;
        RECT 146.715 -28.725 147.045 -28.395 ;
        RECT 142.635 -28.725 142.965 -28.395 ;
        RECT 139.915 -28.725 140.245 -28.395 ;
        RECT 138.555 -28.725 138.885 -28.395 ;
        RECT 134.475 -28.725 134.805 -28.395 ;
        RECT 133.115 -28.725 133.445 -28.395 ;
        RECT 131.755 -28.725 132.085 -28.395 ;
        RECT 127.675 -28.725 128.005 -28.395 ;
        RECT 124.955 -28.725 125.285 -28.395 ;
        RECT 120.875 -28.725 121.205 -28.395 ;
        RECT 119.515 -28.725 119.845 -28.395 ;
        RECT 118.155 -28.725 118.485 -28.395 ;
        RECT 116.795 -28.725 117.125 -28.395 ;
        RECT 112.715 -28.725 113.045 -28.395 ;
        RECT 109.995 -28.725 110.325 -28.395 ;
        RECT 105.915 -28.725 106.245 -28.395 ;
        RECT 104.555 -28.725 104.885 -28.395 ;
        RECT 103.195 -28.725 103.525 -28.395 ;
        RECT 101.835 -28.725 102.165 -28.395 ;
        RECT 97.755 -28.725 98.085 -28.395 ;
        RECT 90.955 -28.725 91.285 -28.395 ;
        RECT 89.595 -28.725 89.925 -28.395 ;
        RECT 88.235 -28.725 88.565 -28.395 ;
        RECT 86.875 -28.725 87.205 -28.395 ;
        RECT 82.795 -28.725 83.125 -28.395 ;
        RECT 80.075 -28.725 80.405 -28.395 ;
        RECT 75.995 -28.725 76.325 -28.395 ;
        RECT 74.635 -28.725 74.965 -28.395 ;
        RECT 73.275 -28.725 73.605 -28.395 ;
        RECT 71.915 -28.725 72.245 -28.395 ;
        RECT 67.835 -28.725 68.165 -28.395 ;
        RECT 65.115 -28.725 65.445 -28.395 ;
        RECT 61.035 -28.725 61.365 -28.395 ;
        RECT 59.675 -28.725 60.005 -28.395 ;
        RECT 58.315 -28.725 58.645 -28.395 ;
        RECT 56.955 -28.725 57.285 -28.395 ;
        RECT 51.515 -28.725 51.845 -28.395 ;
        RECT 50.155 -28.725 50.485 -28.395 ;
        RECT 46.075 -28.725 46.405 -28.395 ;
        RECT 44.715 -28.725 45.045 -28.395 ;
        RECT 43.355 -28.725 43.685 -28.395 ;
        RECT 41.995 -28.725 42.325 -28.395 ;
        RECT 36.555 -28.725 36.885 -28.395 ;
        RECT 35.195 -28.725 35.525 -28.395 ;
        RECT 31.115 -28.725 31.445 -28.395 ;
        RECT 29.755 -28.725 30.085 -28.395 ;
        RECT 28.395 -28.725 28.725 -28.395 ;
        RECT 27.035 -28.725 27.365 -28.395 ;
        RECT 21.595 -28.725 21.925 -28.395 ;
        RECT 20.235 -28.725 20.565 -28.395 ;
        RECT 16.155 -28.725 16.485 -28.395 ;
        RECT 14.795 -28.725 15.125 -28.395 ;
        RECT 13.435 -28.725 13.765 -28.395 ;
        RECT 12.075 -28.725 12.405 -28.395 ;
        RECT 10.715 -28.725 11.045 -28.395 ;
        RECT 7.995 -28.725 8.325 -28.395 ;
        RECT 6.635 -28.725 6.965 -28.395 ;
        RECT 5.275 -28.725 5.605 -28.395 ;
        RECT 3.915 -28.725 4.245 -28.395 ;
        RECT 2.555 -28.725 2.885 -28.395 ;
        RECT 1.195 -28.725 1.525 -28.395 ;
        RECT -0.165 -28.725 0.165 -28.395 ;
        RECT -1.525 -28.725 -1.195 -28.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 954.555 -30.085 954.885 -29.755 ;
        RECT 934.84 -30.08 954.885 -29.76 ;
        RECT 953.195 -30.085 953.525 -29.755 ;
        RECT 951.835 -30.085 952.165 -29.755 ;
        RECT 950.475 -30.085 950.805 -29.755 ;
        RECT 946.395 -30.085 946.725 -29.755 ;
        RECT 945.035 -30.085 945.365 -29.755 ;
        RECT 943.675 -30.085 944.005 -29.755 ;
        RECT 942.315 -30.085 942.645 -29.755 ;
        RECT 940.955 -30.085 941.285 -29.755 ;
        RECT 939.595 -30.085 939.925 -29.755 ;
        RECT 938.235 -30.085 938.565 -29.755 ;
        RECT 936.875 -30.085 937.205 -29.755 ;
        RECT 935.515 -30.085 935.845 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 920.555 -31.445 920.885 -31.115 ;
        RECT 917.835 -31.445 918.165 -31.115 ;
        RECT 915.115 -31.445 915.445 -31.115 ;
        RECT 912.395 -31.445 912.725 -31.115 ;
        RECT 911.035 -31.445 911.365 -31.115 ;
        RECT 909.675 -31.445 910.005 -31.115 ;
        RECT 908.315 -31.445 908.645 -31.115 ;
        RECT 906.955 -31.445 907.285 -31.115 ;
        RECT 905.595 -31.445 905.925 -31.115 ;
        RECT 902.875 -31.445 903.205 -31.115 ;
        RECT 900.155 -31.445 900.485 -31.115 ;
        RECT 897.435 -31.445 897.765 -31.115 ;
        RECT 896.075 -31.445 896.405 -31.115 ;
        RECT 894.715 -31.445 895.045 -31.115 ;
        RECT 893.355 -31.445 893.685 -31.115 ;
        RECT 891.995 -31.445 892.325 -31.115 ;
        RECT 890.635 -31.445 890.965 -31.115 ;
        RECT 887.915 -31.445 888.245 -31.115 ;
        RECT 885.195 -31.445 885.525 -31.115 ;
        RECT 882.475 -31.445 882.805 -31.115 ;
        RECT 881.115 -31.445 881.445 -31.115 ;
        RECT 879.755 -31.445 880.085 -31.115 ;
        RECT 878.395 -31.445 878.725 -31.115 ;
        RECT 877.035 -31.445 877.365 -31.115 ;
        RECT 875.675 -31.445 876.005 -31.115 ;
        RECT 872.955 -31.445 873.285 -31.115 ;
        RECT 870.235 -31.445 870.565 -31.115 ;
        RECT 867.515 -31.445 867.845 -31.115 ;
        RECT 866.155 -31.445 866.485 -31.115 ;
        RECT 864.795 -31.445 865.125 -31.115 ;
        RECT 863.435 -31.445 863.765 -31.115 ;
        RECT 862.075 -31.445 862.405 -31.115 ;
        RECT 860.715 -31.445 861.045 -31.115 ;
        RECT 857.995 -31.445 858.325 -31.115 ;
        RECT 855.275 -31.445 855.605 -31.115 ;
        RECT 852.555 -31.445 852.885 -31.115 ;
        RECT 851.195 -31.445 851.525 -31.115 ;
        RECT 849.835 -31.445 850.165 -31.115 ;
        RECT 848.475 -31.445 848.805 -31.115 ;
        RECT 847.115 -31.445 847.445 -31.115 ;
        RECT 845.755 -31.445 846.085 -31.115 ;
        RECT 843.035 -31.445 843.365 -31.115 ;
        RECT 840.315 -31.445 840.645 -31.115 ;
        RECT 837.595 -31.445 837.925 -31.115 ;
        RECT 836.235 -31.445 836.565 -31.115 ;
        RECT 834.875 -31.445 835.205 -31.115 ;
        RECT 833.515 -31.445 833.845 -31.115 ;
        RECT 832.155 -31.445 832.485 -31.115 ;
        RECT 828.075 -31.445 828.405 -31.115 ;
        RECT 825.355 -31.445 825.685 -31.115 ;
        RECT 822.635 -31.445 822.965 -31.115 ;
        RECT 821.275 -31.445 821.605 -31.115 ;
        RECT 819.915 -31.445 820.245 -31.115 ;
        RECT 818.555 -31.445 818.885 -31.115 ;
        RECT 817.195 -31.445 817.525 -31.115 ;
        RECT 813.115 -31.445 813.445 -31.115 ;
        RECT 810.395 -31.445 810.725 -31.115 ;
        RECT 807.675 -31.445 808.005 -31.115 ;
        RECT 806.315 -31.445 806.645 -31.115 ;
        RECT 804.955 -31.445 805.285 -31.115 ;
        RECT 803.595 -31.445 803.925 -31.115 ;
        RECT 802.235 -31.445 802.565 -31.115 ;
        RECT 798.155 -31.445 798.485 -31.115 ;
        RECT 795.435 -31.445 795.765 -31.115 ;
        RECT 792.715 -31.445 793.045 -31.115 ;
        RECT 791.355 -31.445 791.685 -31.115 ;
        RECT 789.995 -31.445 790.325 -31.115 ;
        RECT 788.635 -31.445 788.965 -31.115 ;
        RECT 787.275 -31.445 787.605 -31.115 ;
        RECT 783.195 -31.445 783.525 -31.115 ;
        RECT 780.475 -31.445 780.805 -31.115 ;
        RECT 779.115 -31.445 779.445 -31.115 ;
        RECT 777.755 -31.445 778.085 -31.115 ;
        RECT 776.395 -31.445 776.725 -31.115 ;
        RECT 775.035 -31.445 775.365 -31.115 ;
        RECT 773.675 -31.445 774.005 -31.115 ;
        RECT 772.315 -31.445 772.645 -31.115 ;
        RECT 768.235 -31.445 768.565 -31.115 ;
        RECT 764.155 -31.445 764.485 -31.115 ;
        RECT 762.795 -31.445 763.125 -31.115 ;
        RECT 761.435 -31.445 761.765 -31.115 ;
        RECT 760.075 -31.445 760.405 -31.115 ;
        RECT 758.715 -31.445 759.045 -31.115 ;
        RECT 757.355 -31.445 757.685 -31.115 ;
        RECT 753.275 -31.445 753.605 -31.115 ;
        RECT 749.195 -31.445 749.525 -31.115 ;
        RECT 747.835 -31.445 748.165 -31.115 ;
        RECT 746.475 -31.445 746.805 -31.115 ;
        RECT 745.115 -31.445 745.445 -31.115 ;
        RECT 743.755 -31.445 744.085 -31.115 ;
        RECT 742.395 -31.445 742.725 -31.115 ;
        RECT 738.315 -31.445 738.645 -31.115 ;
        RECT 734.235 -31.445 734.565 -31.115 ;
        RECT 732.875 -31.445 733.205 -31.115 ;
        RECT 731.515 -31.445 731.845 -31.115 ;
        RECT 730.155 -31.445 730.485 -31.115 ;
        RECT 728.795 -31.445 729.125 -31.115 ;
        RECT 727.435 -31.445 727.765 -31.115 ;
        RECT 721.995 -31.445 722.325 -31.115 ;
        RECT 719.275 -31.445 719.605 -31.115 ;
        RECT 717.915 -31.445 718.245 -31.115 ;
        RECT 716.555 -31.445 716.885 -31.115 ;
        RECT 715.195 -31.445 715.525 -31.115 ;
        RECT 713.835 -31.445 714.165 -31.115 ;
        RECT 712.475 -31.445 712.805 -31.115 ;
        RECT 707.035 -31.445 707.365 -31.115 ;
        RECT 704.315 -31.445 704.645 -31.115 ;
        RECT 702.955 -31.445 703.285 -31.115 ;
        RECT 701.595 -31.445 701.925 -31.115 ;
        RECT 700.235 -31.445 700.565 -31.115 ;
        RECT 698.875 -31.445 699.205 -31.115 ;
        RECT 697.515 -31.445 697.845 -31.115 ;
        RECT 692.075 -31.445 692.405 -31.115 ;
        RECT 689.355 -31.445 689.685 -31.115 ;
        RECT 687.995 -31.445 688.325 -31.115 ;
        RECT 686.635 -31.445 686.965 -31.115 ;
        RECT 685.275 -31.445 685.605 -31.115 ;
        RECT 683.915 -31.445 684.245 -31.115 ;
        RECT 682.555 -31.445 682.885 -31.115 ;
        RECT 679.835 -31.445 680.165 -31.115 ;
        RECT 677.115 -31.445 677.445 -31.115 ;
        RECT 674.395 -31.445 674.725 -31.115 ;
        RECT 673.035 -31.445 673.365 -31.115 ;
        RECT 671.675 -31.445 672.005 -31.115 ;
        RECT 670.315 -31.445 670.645 -31.115 ;
        RECT 668.955 -31.445 669.285 -31.115 ;
        RECT 667.595 -31.445 667.925 -31.115 ;
        RECT 664.875 -31.445 665.205 -31.115 ;
        RECT 662.155 -31.445 662.485 -31.115 ;
        RECT 659.435 -31.445 659.765 -31.115 ;
        RECT 658.075 -31.445 658.405 -31.115 ;
        RECT 656.715 -31.445 657.045 -31.115 ;
        RECT 655.355 -31.445 655.685 -31.115 ;
        RECT 653.995 -31.445 654.325 -31.115 ;
        RECT 652.635 -31.445 652.965 -31.115 ;
        RECT 649.915 -31.445 650.245 -31.115 ;
        RECT 647.195 -31.445 647.525 -31.115 ;
        RECT 644.475 -31.445 644.805 -31.115 ;
        RECT 643.115 -31.445 643.445 -31.115 ;
        RECT 641.755 -31.445 642.085 -31.115 ;
        RECT 640.395 -31.445 640.725 -31.115 ;
        RECT 639.035 -31.445 639.365 -31.115 ;
        RECT 637.675 -31.445 638.005 -31.115 ;
        RECT 634.955 -31.445 635.285 -31.115 ;
        RECT 632.235 -31.445 632.565 -31.115 ;
        RECT 629.515 -31.445 629.845 -31.115 ;
        RECT 628.155 -31.445 628.485 -31.115 ;
        RECT 626.795 -31.445 627.125 -31.115 ;
        RECT 625.435 -31.445 625.765 -31.115 ;
        RECT 624.075 -31.445 624.405 -31.115 ;
        RECT 622.715 -31.445 623.045 -31.115 ;
        RECT 619.995 -31.445 620.325 -31.115 ;
        RECT 617.275 -31.445 617.605 -31.115 ;
        RECT 614.555 -31.445 614.885 -31.115 ;
        RECT 613.195 -31.445 613.525 -31.115 ;
        RECT 611.835 -31.445 612.165 -31.115 ;
        RECT 610.475 -31.445 610.805 -31.115 ;
        RECT 609.115 -31.445 609.445 -31.115 ;
        RECT 607.755 -31.445 608.085 -31.115 ;
        RECT 605.035 -31.445 605.365 -31.115 ;
        RECT 602.315 -31.445 602.645 -31.115 ;
        RECT 599.595 -31.445 599.925 -31.115 ;
        RECT 598.235 -31.445 598.565 -31.115 ;
        RECT 596.875 -31.445 597.205 -31.115 ;
        RECT 595.515 -31.445 595.845 -31.115 ;
        RECT 594.155 -31.445 594.485 -31.115 ;
        RECT 592.795 -31.445 593.125 -31.115 ;
        RECT 590.075 -31.445 590.405 -31.115 ;
        RECT 587.355 -31.445 587.685 -31.115 ;
        RECT 584.635 -31.445 584.965 -31.115 ;
        RECT 583.275 -31.445 583.605 -31.115 ;
        RECT 581.915 -31.445 582.245 -31.115 ;
        RECT 580.555 -31.445 580.885 -31.115 ;
        RECT 579.195 -31.445 579.525 -31.115 ;
        RECT 577.835 -31.445 578.165 -31.115 ;
        RECT 575.115 -31.445 575.445 -31.115 ;
        RECT 572.395 -31.445 572.725 -31.115 ;
        RECT 569.675 -31.445 570.005 -31.115 ;
        RECT 568.315 -31.445 568.645 -31.115 ;
        RECT 566.955 -31.445 567.285 -31.115 ;
        RECT 565.595 -31.445 565.925 -31.115 ;
        RECT 564.235 -31.445 564.565 -31.115 ;
        RECT 562.875 -31.445 563.205 -31.115 ;
        RECT 560.155 -31.445 560.485 -31.115 ;
        RECT 557.435 -31.445 557.765 -31.115 ;
        RECT 554.715 -31.445 555.045 -31.115 ;
        RECT 553.355 -31.445 553.685 -31.115 ;
        RECT 551.995 -31.445 552.325 -31.115 ;
        RECT 550.635 -31.445 550.965 -31.115 ;
        RECT 549.275 -31.445 549.605 -31.115 ;
        RECT 547.915 -31.445 548.245 -31.115 ;
        RECT 545.195 -31.445 545.525 -31.115 ;
        RECT 542.475 -31.445 542.805 -31.115 ;
        RECT 539.755 -31.445 540.085 -31.115 ;
        RECT 538.395 -31.445 538.725 -31.115 ;
        RECT 537.035 -31.445 537.365 -31.115 ;
        RECT 535.675 -31.445 536.005 -31.115 ;
        RECT 534.315 -31.445 534.645 -31.115 ;
        RECT 532.955 -31.445 533.285 -31.115 ;
        RECT 530.235 -31.445 530.565 -31.115 ;
        RECT 527.515 -31.445 527.845 -31.115 ;
        RECT 524.795 -31.445 525.125 -31.115 ;
        RECT 523.435 -31.445 523.765 -31.115 ;
        RECT 522.075 -31.445 522.405 -31.115 ;
        RECT 520.715 -31.445 521.045 -31.115 ;
        RECT 519.355 -31.445 519.685 -31.115 ;
        RECT 517.995 -31.445 518.325 -31.115 ;
        RECT 515.275 -31.445 515.605 -31.115 ;
        RECT 512.555 -31.445 512.885 -31.115 ;
        RECT 509.835 -31.445 510.165 -31.115 ;
        RECT 508.475 -31.445 508.805 -31.115 ;
        RECT 507.115 -31.445 507.445 -31.115 ;
        RECT 505.755 -31.445 506.085 -31.115 ;
        RECT 504.395 -31.445 504.725 -31.115 ;
        RECT 500.315 -31.445 500.645 -31.115 ;
        RECT 497.595 -31.445 497.925 -31.115 ;
        RECT 494.875 -31.445 495.205 -31.115 ;
        RECT 493.515 -31.445 493.845 -31.115 ;
        RECT 492.155 -31.445 492.485 -31.115 ;
        RECT 490.795 -31.445 491.125 -31.115 ;
        RECT 489.435 -31.445 489.765 -31.115 ;
        RECT 485.355 -31.445 485.685 -31.115 ;
        RECT 482.635 -31.445 482.965 -31.115 ;
        RECT 479.915 -31.445 480.245 -31.115 ;
        RECT 478.555 -31.445 478.885 -31.115 ;
        RECT 477.195 -31.445 477.525 -31.115 ;
        RECT 475.835 -31.445 476.165 -31.115 ;
        RECT 474.475 -31.445 474.805 -31.115 ;
        RECT 470.395 -31.445 470.725 -31.115 ;
        RECT 467.675 -31.445 468.005 -31.115 ;
        RECT 464.955 -31.445 465.285 -31.115 ;
        RECT 463.595 -31.445 463.925 -31.115 ;
        RECT 462.235 -31.445 462.565 -31.115 ;
        RECT 460.875 -31.445 461.205 -31.115 ;
        RECT 459.515 -31.445 459.845 -31.115 ;
        RECT 455.435 -31.445 455.765 -31.115 ;
        RECT 452.715 -31.445 453.045 -31.115 ;
        RECT 449.995 -31.445 450.325 -31.115 ;
        RECT 448.635 -31.445 448.965 -31.115 ;
        RECT 447.275 -31.445 447.605 -31.115 ;
        RECT 445.915 -31.445 446.245 -31.115 ;
        RECT 444.555 -31.445 444.885 -31.115 ;
        RECT 440.475 -31.445 440.805 -31.115 ;
        RECT 436.395 -31.445 436.725 -31.115 ;
        RECT 435.035 -31.445 435.365 -31.115 ;
        RECT 433.675 -31.445 434.005 -31.115 ;
        RECT 432.315 -31.445 432.645 -31.115 ;
        RECT 430.955 -31.445 431.285 -31.115 ;
        RECT 429.595 -31.445 429.925 -31.115 ;
        RECT 425.515 -31.445 425.845 -31.115 ;
        RECT 421.435 -31.445 421.765 -31.115 ;
        RECT 420.075 -31.445 420.405 -31.115 ;
        RECT 418.715 -31.445 419.045 -31.115 ;
        RECT 417.355 -31.445 417.685 -31.115 ;
        RECT 415.995 -31.445 416.325 -31.115 ;
        RECT 414.635 -31.445 414.965 -31.115 ;
        RECT 410.555 -31.445 410.885 -31.115 ;
        RECT 406.475 -31.445 406.805 -31.115 ;
        RECT 405.115 -31.445 405.445 -31.115 ;
        RECT 403.755 -31.445 404.085 -31.115 ;
        RECT 402.395 -31.445 402.725 -31.115 ;
        RECT 401.035 -31.445 401.365 -31.115 ;
        RECT 399.675 -31.445 400.005 -31.115 ;
        RECT 395.595 -31.445 395.925 -31.115 ;
        RECT 394.235 -31.445 394.565 -31.115 ;
        RECT 391.515 -31.445 391.845 -31.115 ;
        RECT 390.155 -31.445 390.485 -31.115 ;
        RECT 388.795 -31.445 389.125 -31.115 ;
        RECT 387.435 -31.445 387.765 -31.115 ;
        RECT 386.075 -31.445 386.405 -31.115 ;
        RECT 384.715 -31.445 385.045 -31.115 ;
        RECT 379.275 -31.445 379.605 -31.115 ;
        RECT 376.555 -31.445 376.885 -31.115 ;
        RECT 375.195 -31.445 375.525 -31.115 ;
        RECT 373.835 -31.445 374.165 -31.115 ;
        RECT 372.475 -31.445 372.805 -31.115 ;
        RECT 371.115 -31.445 371.445 -31.115 ;
        RECT 369.755 -31.445 370.085 -31.115 ;
        RECT 364.315 -31.445 364.645 -31.115 ;
        RECT 361.595 -31.445 361.925 -31.115 ;
        RECT 360.235 -31.445 360.565 -31.115 ;
        RECT 358.875 -31.445 359.205 -31.115 ;
        RECT 357.515 -31.445 357.845 -31.115 ;
        RECT 356.155 -31.445 356.485 -31.115 ;
        RECT 354.795 -31.445 355.125 -31.115 ;
        RECT 349.355 -31.445 349.685 -31.115 ;
        RECT 346.635 -31.445 346.965 -31.115 ;
        RECT 345.275 -31.445 345.605 -31.115 ;
        RECT 343.915 -31.445 344.245 -31.115 ;
        RECT 342.555 -31.445 342.885 -31.115 ;
        RECT 341.195 -31.445 341.525 -31.115 ;
        RECT 339.835 -31.445 340.165 -31.115 ;
        RECT 337.115 -31.445 337.445 -31.115 ;
        RECT 334.395 -31.445 334.725 -31.115 ;
        RECT 331.675 -31.445 332.005 -31.115 ;
        RECT 330.315 -31.445 330.645 -31.115 ;
        RECT 328.955 -31.445 329.285 -31.115 ;
        RECT 327.595 -31.445 327.925 -31.115 ;
        RECT 326.235 -31.445 326.565 -31.115 ;
        RECT 324.875 -31.445 325.205 -31.115 ;
        RECT 322.155 -31.445 322.485 -31.115 ;
        RECT 319.435 -31.445 319.765 -31.115 ;
        RECT 316.715 -31.445 317.045 -31.115 ;
        RECT 315.355 -31.445 315.685 -31.115 ;
        RECT 313.995 -31.445 314.325 -31.115 ;
        RECT 312.635 -31.445 312.965 -31.115 ;
        RECT 311.275 -31.445 311.605 -31.115 ;
        RECT 309.915 -31.445 310.245 -31.115 ;
        RECT 307.195 -31.445 307.525 -31.115 ;
        RECT 304.475 -31.445 304.805 -31.115 ;
        RECT 301.755 -31.445 302.085 -31.115 ;
        RECT 300.395 -31.445 300.725 -31.115 ;
        RECT 299.035 -31.445 299.365 -31.115 ;
        RECT 297.675 -31.445 298.005 -31.115 ;
        RECT 296.315 -31.445 296.645 -31.115 ;
        RECT 294.955 -31.445 295.285 -31.115 ;
        RECT 292.235 -31.445 292.565 -31.115 ;
        RECT 289.515 -31.445 289.845 -31.115 ;
        RECT 286.795 -31.445 287.125 -31.115 ;
        RECT 285.435 -31.445 285.765 -31.115 ;
        RECT 284.075 -31.445 284.405 -31.115 ;
        RECT 282.715 -31.445 283.045 -31.115 ;
        RECT 281.355 -31.445 281.685 -31.115 ;
        RECT 279.995 -31.445 280.325 -31.115 ;
        RECT 277.275 -31.445 277.605 -31.115 ;
        RECT 274.555 -31.445 274.885 -31.115 ;
        RECT 271.835 -31.445 272.165 -31.115 ;
        RECT 270.475 -31.445 270.805 -31.115 ;
        RECT 269.115 -31.445 269.445 -31.115 ;
        RECT 267.755 -31.445 268.085 -31.115 ;
        RECT 266.395 -31.445 266.725 -31.115 ;
        RECT 265.035 -31.445 265.365 -31.115 ;
        RECT 262.315 -31.445 262.645 -31.115 ;
        RECT 259.595 -31.445 259.925 -31.115 ;
        RECT 256.875 -31.445 257.205 -31.115 ;
        RECT 255.515 -31.445 255.845 -31.115 ;
        RECT 254.155 -31.445 254.485 -31.115 ;
        RECT 252.795 -31.445 253.125 -31.115 ;
        RECT 251.435 -31.445 251.765 -31.115 ;
        RECT 250.075 -31.445 250.405 -31.115 ;
        RECT 247.355 -31.445 247.685 -31.115 ;
        RECT 244.635 -31.445 244.965 -31.115 ;
        RECT 241.915 -31.445 242.245 -31.115 ;
        RECT 240.555 -31.445 240.885 -31.115 ;
        RECT 239.195 -31.445 239.525 -31.115 ;
        RECT 237.835 -31.445 238.165 -31.115 ;
        RECT 236.475 -31.445 236.805 -31.115 ;
        RECT 235.115 -31.445 235.445 -31.115 ;
        RECT 232.395 -31.445 232.725 -31.115 ;
        RECT 229.675 -31.445 230.005 -31.115 ;
        RECT 226.955 -31.445 227.285 -31.115 ;
        RECT 225.595 -31.445 225.925 -31.115 ;
        RECT 224.235 -31.445 224.565 -31.115 ;
        RECT 222.875 -31.445 223.205 -31.115 ;
        RECT 221.515 -31.445 221.845 -31.115 ;
        RECT 220.155 -31.445 220.485 -31.115 ;
        RECT 217.435 -31.445 217.765 -31.115 ;
        RECT 214.715 -31.445 215.045 -31.115 ;
        RECT 211.995 -31.445 212.325 -31.115 ;
        RECT 210.635 -31.445 210.965 -31.115 ;
        RECT 209.275 -31.445 209.605 -31.115 ;
        RECT 207.915 -31.445 208.245 -31.115 ;
        RECT 206.555 -31.445 206.885 -31.115 ;
        RECT 205.195 -31.445 205.525 -31.115 ;
        RECT 202.475 -31.445 202.805 -31.115 ;
        RECT 199.755 -31.445 200.085 -31.115 ;
        RECT 197.035 -31.445 197.365 -31.115 ;
        RECT 195.675 -31.445 196.005 -31.115 ;
        RECT 194.315 -31.445 194.645 -31.115 ;
        RECT 192.955 -31.445 193.285 -31.115 ;
        RECT 191.595 -31.445 191.925 -31.115 ;
        RECT 190.235 -31.445 190.565 -31.115 ;
        RECT 187.515 -31.445 187.845 -31.115 ;
        RECT 184.795 -31.445 185.125 -31.115 ;
        RECT 182.075 -31.445 182.405 -31.115 ;
        RECT 180.715 -31.445 181.045 -31.115 ;
        RECT 179.355 -31.445 179.685 -31.115 ;
        RECT 177.995 -31.445 178.325 -31.115 ;
        RECT 176.635 -31.445 176.965 -31.115 ;
        RECT 175.275 -31.445 175.605 -31.115 ;
        RECT 172.555 -31.445 172.885 -31.115 ;
        RECT 169.835 -31.445 170.165 -31.115 ;
        RECT 167.115 -31.445 167.445 -31.115 ;
        RECT 165.755 -31.445 166.085 -31.115 ;
        RECT 164.395 -31.445 164.725 -31.115 ;
        RECT 163.035 -31.445 163.365 -31.115 ;
        RECT 161.675 -31.445 162.005 -31.115 ;
        RECT 157.595 -31.445 157.925 -31.115 ;
        RECT 154.875 -31.445 155.205 -31.115 ;
        RECT 152.155 -31.445 152.485 -31.115 ;
        RECT 150.795 -31.445 151.125 -31.115 ;
        RECT 149.435 -31.445 149.765 -31.115 ;
        RECT 148.075 -31.445 148.405 -31.115 ;
        RECT 146.715 -31.445 147.045 -31.115 ;
        RECT 142.635 -31.445 142.965 -31.115 ;
        RECT 139.915 -31.445 140.245 -31.115 ;
        RECT 137.195 -31.445 137.525 -31.115 ;
        RECT 135.835 -31.445 136.165 -31.115 ;
        RECT 134.475 -31.445 134.805 -31.115 ;
        RECT 133.115 -31.445 133.445 -31.115 ;
        RECT 131.755 -31.445 132.085 -31.115 ;
        RECT 127.675 -31.445 128.005 -31.115 ;
        RECT 124.955 -31.445 125.285 -31.115 ;
        RECT 122.235 -31.445 122.565 -31.115 ;
        RECT 120.875 -31.445 121.205 -31.115 ;
        RECT 119.515 -31.445 119.845 -31.115 ;
        RECT 118.155 -31.445 118.485 -31.115 ;
        RECT 116.795 -31.445 117.125 -31.115 ;
        RECT 112.715 -31.445 113.045 -31.115 ;
        RECT 109.995 -31.445 110.325 -31.115 ;
        RECT 107.275 -31.445 107.605 -31.115 ;
        RECT 105.915 -31.445 106.245 -31.115 ;
        RECT 104.555 -31.445 104.885 -31.115 ;
        RECT 103.195 -31.445 103.525 -31.115 ;
        RECT 101.835 -31.445 102.165 -31.115 ;
        RECT 97.755 -31.445 98.085 -31.115 ;
        RECT 93.675 -31.445 94.005 -31.115 ;
        RECT 92.315 -31.445 92.645 -31.115 ;
        RECT 90.955 -31.445 91.285 -31.115 ;
        RECT 89.595 -31.445 89.925 -31.115 ;
        RECT 88.235 -31.445 88.565 -31.115 ;
        RECT 86.875 -31.445 87.205 -31.115 ;
        RECT 82.795 -31.445 83.125 -31.115 ;
        RECT 78.715 -31.445 79.045 -31.115 ;
        RECT 77.355 -31.445 77.685 -31.115 ;
        RECT 75.995 -31.445 76.325 -31.115 ;
        RECT 74.635 -31.445 74.965 -31.115 ;
        RECT 73.275 -31.445 73.605 -31.115 ;
        RECT 71.915 -31.445 72.245 -31.115 ;
        RECT 67.835 -31.445 68.165 -31.115 ;
        RECT 63.755 -31.445 64.085 -31.115 ;
        RECT 62.395 -31.445 62.725 -31.115 ;
        RECT 61.035 -31.445 61.365 -31.115 ;
        RECT 59.675 -31.445 60.005 -31.115 ;
        RECT 58.315 -31.445 58.645 -31.115 ;
        RECT 56.955 -31.445 57.285 -31.115 ;
        RECT 51.515 -31.445 51.845 -31.115 ;
        RECT 48.795 -31.445 49.125 -31.115 ;
        RECT 47.435 -31.445 47.765 -31.115 ;
        RECT 46.075 -31.445 46.405 -31.115 ;
        RECT 44.715 -31.445 45.045 -31.115 ;
        RECT 43.355 -31.445 43.685 -31.115 ;
        RECT 41.995 -31.445 42.325 -31.115 ;
        RECT 36.555 -31.445 36.885 -31.115 ;
        RECT 33.835 -31.445 34.165 -31.115 ;
        RECT 32.475 -31.445 32.805 -31.115 ;
        RECT 31.115 -31.445 31.445 -31.115 ;
        RECT 29.755 -31.445 30.085 -31.115 ;
        RECT 28.395 -31.445 28.725 -31.115 ;
        RECT 27.035 -31.445 27.365 -31.115 ;
        RECT 21.595 -31.445 21.925 -31.115 ;
        RECT 18.875 -31.445 19.205 -31.115 ;
        RECT 17.515 -31.445 17.845 -31.115 ;
        RECT 16.155 -31.445 16.485 -31.115 ;
        RECT 14.795 -31.445 15.125 -31.115 ;
        RECT 13.435 -31.445 13.765 -31.115 ;
        RECT 12.075 -31.445 12.405 -31.115 ;
        RECT 10.715 -31.445 11.045 -31.115 ;
        RECT 7.995 -31.445 8.325 -31.115 ;
        RECT 6.635 -31.445 6.965 -31.115 ;
        RECT 5.275 -31.445 5.605 -31.115 ;
        RECT 3.915 -31.445 4.245 -31.115 ;
        RECT 2.555 -31.445 2.885 -31.115 ;
        RECT 1.195 -31.445 1.525 -31.115 ;
        RECT -0.165 -31.445 0.165 -31.115 ;
        RECT -1.525 -31.445 -1.195 -31.115 ;
        RECT 954.555 -31.445 954.885 -31.115 ;
        RECT -1.525 -31.44 954.885 -31.12 ;
        RECT 953.195 -31.445 953.525 -31.115 ;
        RECT 951.835 -31.445 952.165 -31.115 ;
        RECT 950.475 -31.445 950.805 -31.115 ;
        RECT 946.395 -31.445 946.725 -31.115 ;
        RECT 945.035 -31.445 945.365 -31.115 ;
        RECT 943.675 -31.445 944.005 -31.115 ;
        RECT 942.315 -31.445 942.645 -31.115 ;
        RECT 940.955 -31.445 941.285 -31.115 ;
        RECT 939.595 -31.445 939.925 -31.115 ;
        RECT 938.235 -31.445 938.565 -31.115 ;
        RECT 936.875 -31.445 937.205 -31.115 ;
        RECT 935.515 -31.445 935.845 -31.115 ;
        RECT 932.795 -31.445 933.125 -31.115 ;
        RECT 930.075 -31.445 930.405 -31.115 ;
        RECT 927.355 -31.445 927.685 -31.115 ;
        RECT 925.995 -31.445 926.325 -31.115 ;
        RECT 924.635 -31.445 924.965 -31.115 ;
        RECT 923.275 -31.445 923.605 -31.115 ;
        RECT 921.915 -31.445 922.245 -31.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 916.48 -27.36 927 -27.04 ;
        RECT 924.635 -27.365 924.965 -27.035 ;
        RECT 923.275 -27.365 923.605 -27.035 ;
        RECT 921.915 -27.365 922.245 -27.035 ;
        RECT 920.555 -27.365 920.885 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 919.88 -35.52 927 -35.2 ;
        RECT 925.995 -35.525 926.325 -35.195 ;
        RECT 924.635 -35.525 924.965 -35.195 ;
        RECT 923.275 -35.525 923.605 -35.195 ;
        RECT 921.915 -35.525 922.245 -35.195 ;
        RECT 920.555 -35.525 920.885 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 919.88 -26 930.4 -25.68 ;
        RECT 928.715 -26.005 929.045 -25.675 ;
        RECT 924.635 -26.005 924.965 -25.675 ;
        RECT 923.275 -26.005 923.605 -25.675 ;
        RECT 921.915 -26.005 922.245 -25.675 ;
        RECT 920.555 -26.005 920.885 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 930.76 -23.28 941.28 -22.96 ;
        RECT 939.595 -23.285 939.925 -22.955 ;
        RECT 938.235 -23.285 938.565 -22.955 ;
        RECT 936.875 -23.285 937.205 -22.955 ;
        RECT 935.515 -23.285 935.845 -22.955 ;
        RECT 931.435 -23.285 931.765 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 943.675 -35.525 944.005 -35.195 ;
        RECT 934.84 -35.52 944.005 -35.2 ;
        RECT 942.315 -35.525 942.645 -35.195 ;
        RECT 940.955 -35.525 941.285 -35.195 ;
        RECT 939.595 -35.525 939.925 -35.195 ;
        RECT 938.235 -35.525 938.565 -35.195 ;
        RECT 936.875 -35.525 937.205 -35.195 ;
        RECT 935.515 -35.525 935.845 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -20.56 920.555 -20.24 ;
        RECT 919.195 -20.565 919.525 -20.235 ;
        RECT 917.835 -20.565 918.165 -20.235 ;
        RECT 916.475 -20.565 916.805 -20.235 ;
        RECT 911.035 -20.565 911.365 -20.235 ;
        RECT 909.675 -20.565 910.005 -20.235 ;
        RECT 908.315 -20.565 908.645 -20.235 ;
        RECT 906.955 -20.565 907.285 -20.235 ;
        RECT 905.595 -20.565 905.925 -20.235 ;
        RECT 904.235 -20.565 904.565 -20.235 ;
        RECT 902.875 -20.565 903.205 -20.235 ;
        RECT 901.515 -20.565 901.845 -20.235 ;
        RECT 896.075 -20.565 896.405 -20.235 ;
        RECT 894.715 -20.565 895.045 -20.235 ;
        RECT 893.355 -20.565 893.685 -20.235 ;
        RECT 891.995 -20.565 892.325 -20.235 ;
        RECT 890.635 -20.565 890.965 -20.235 ;
        RECT 889.275 -20.565 889.605 -20.235 ;
        RECT 887.915 -20.565 888.245 -20.235 ;
        RECT 886.555 -20.565 886.885 -20.235 ;
        RECT 881.115 -20.565 881.445 -20.235 ;
        RECT 879.755 -20.565 880.085 -20.235 ;
        RECT 878.395 -20.565 878.725 -20.235 ;
        RECT 877.035 -20.565 877.365 -20.235 ;
        RECT 875.675 -20.565 876.005 -20.235 ;
        RECT 874.315 -20.565 874.645 -20.235 ;
        RECT 872.955 -20.565 873.285 -20.235 ;
        RECT 871.595 -20.565 871.925 -20.235 ;
        RECT 866.155 -20.565 866.485 -20.235 ;
        RECT 864.795 -20.565 865.125 -20.235 ;
        RECT 863.435 -20.565 863.765 -20.235 ;
        RECT 862.075 -20.565 862.405 -20.235 ;
        RECT 860.715 -20.565 861.045 -20.235 ;
        RECT 859.355 -20.565 859.685 -20.235 ;
        RECT 857.995 -20.565 858.325 -20.235 ;
        RECT 856.635 -20.565 856.965 -20.235 ;
        RECT 851.195 -20.565 851.525 -20.235 ;
        RECT 849.835 -20.565 850.165 -20.235 ;
        RECT 848.475 -20.565 848.805 -20.235 ;
        RECT 847.115 -20.565 847.445 -20.235 ;
        RECT 845.755 -20.565 846.085 -20.235 ;
        RECT 844.395 -20.565 844.725 -20.235 ;
        RECT 843.035 -20.565 843.365 -20.235 ;
        RECT 841.675 -20.565 842.005 -20.235 ;
        RECT 836.235 -20.565 836.565 -20.235 ;
        RECT 834.875 -20.565 835.205 -20.235 ;
        RECT 833.515 -20.565 833.845 -20.235 ;
        RECT 832.155 -20.565 832.485 -20.235 ;
        RECT 830.795 -20.565 831.125 -20.235 ;
        RECT 829.435 -20.565 829.765 -20.235 ;
        RECT 828.075 -20.565 828.405 -20.235 ;
        RECT 826.715 -20.565 827.045 -20.235 ;
        RECT 821.275 -20.565 821.605 -20.235 ;
        RECT 819.915 -20.565 820.245 -20.235 ;
        RECT 818.555 -20.565 818.885 -20.235 ;
        RECT 817.195 -20.565 817.525 -20.235 ;
        RECT 815.835 -20.565 816.165 -20.235 ;
        RECT 814.475 -20.565 814.805 -20.235 ;
        RECT 813.115 -20.565 813.445 -20.235 ;
        RECT 811.755 -20.565 812.085 -20.235 ;
        RECT 806.315 -20.565 806.645 -20.235 ;
        RECT 804.955 -20.565 805.285 -20.235 ;
        RECT 803.595 -20.565 803.925 -20.235 ;
        RECT 802.235 -20.565 802.565 -20.235 ;
        RECT 800.875 -20.565 801.205 -20.235 ;
        RECT 799.515 -20.565 799.845 -20.235 ;
        RECT 798.155 -20.565 798.485 -20.235 ;
        RECT 796.795 -20.565 797.125 -20.235 ;
        RECT 791.355 -20.565 791.685 -20.235 ;
        RECT 789.995 -20.565 790.325 -20.235 ;
        RECT 788.635 -20.565 788.965 -20.235 ;
        RECT 787.275 -20.565 787.605 -20.235 ;
        RECT 785.915 -20.565 786.245 -20.235 ;
        RECT 784.555 -20.565 784.885 -20.235 ;
        RECT 783.195 -20.565 783.525 -20.235 ;
        RECT 781.835 -20.565 782.165 -20.235 ;
        RECT 779.115 -20.565 779.445 -20.235 ;
        RECT 776.395 -20.565 776.725 -20.235 ;
        RECT 775.035 -20.565 775.365 -20.235 ;
        RECT 773.675 -20.565 774.005 -20.235 ;
        RECT 772.315 -20.565 772.645 -20.235 ;
        RECT 770.955 -20.565 771.285 -20.235 ;
        RECT 769.595 -20.565 769.925 -20.235 ;
        RECT 768.235 -20.565 768.565 -20.235 ;
        RECT 766.875 -20.565 767.205 -20.235 ;
        RECT 764.155 -20.565 764.485 -20.235 ;
        RECT 761.435 -20.565 761.765 -20.235 ;
        RECT 760.075 -20.565 760.405 -20.235 ;
        RECT 758.715 -20.565 759.045 -20.235 ;
        RECT 757.355 -20.565 757.685 -20.235 ;
        RECT 755.995 -20.565 756.325 -20.235 ;
        RECT 754.635 -20.565 754.965 -20.235 ;
        RECT 753.275 -20.565 753.605 -20.235 ;
        RECT 749.195 -20.565 749.525 -20.235 ;
        RECT 746.475 -20.565 746.805 -20.235 ;
        RECT 745.115 -20.565 745.445 -20.235 ;
        RECT 743.755 -20.565 744.085 -20.235 ;
        RECT 742.395 -20.565 742.725 -20.235 ;
        RECT 741.035 -20.565 741.365 -20.235 ;
        RECT 739.675 -20.565 740.005 -20.235 ;
        RECT 738.315 -20.565 738.645 -20.235 ;
        RECT 734.235 -20.565 734.565 -20.235 ;
        RECT 731.515 -20.565 731.845 -20.235 ;
        RECT 730.155 -20.565 730.485 -20.235 ;
        RECT 728.795 -20.565 729.125 -20.235 ;
        RECT 727.435 -20.565 727.765 -20.235 ;
        RECT 726.075 -20.565 726.405 -20.235 ;
        RECT 724.715 -20.565 725.045 -20.235 ;
        RECT 723.355 -20.565 723.685 -20.235 ;
        RECT 719.275 -20.565 719.605 -20.235 ;
        RECT 716.555 -20.565 716.885 -20.235 ;
        RECT 715.195 -20.565 715.525 -20.235 ;
        RECT 713.835 -20.565 714.165 -20.235 ;
        RECT 712.475 -20.565 712.805 -20.235 ;
        RECT 711.115 -20.565 711.445 -20.235 ;
        RECT 709.755 -20.565 710.085 -20.235 ;
        RECT 708.395 -20.565 708.725 -20.235 ;
        RECT 704.315 -20.565 704.645 -20.235 ;
        RECT 701.595 -20.565 701.925 -20.235 ;
        RECT 700.235 -20.565 700.565 -20.235 ;
        RECT 698.875 -20.565 699.205 -20.235 ;
        RECT 697.515 -20.565 697.845 -20.235 ;
        RECT 696.155 -20.565 696.485 -20.235 ;
        RECT 694.795 -20.565 695.125 -20.235 ;
        RECT 693.435 -20.565 693.765 -20.235 ;
        RECT 689.355 -20.565 689.685 -20.235 ;
        RECT 686.635 -20.565 686.965 -20.235 ;
        RECT 685.275 -20.565 685.605 -20.235 ;
        RECT 683.915 -20.565 684.245 -20.235 ;
        RECT 682.555 -20.565 682.885 -20.235 ;
        RECT 681.195 -20.565 681.525 -20.235 ;
        RECT 679.835 -20.565 680.165 -20.235 ;
        RECT 678.475 -20.565 678.805 -20.235 ;
        RECT 674.395 -20.565 674.725 -20.235 ;
        RECT 671.675 -20.565 672.005 -20.235 ;
        RECT 670.315 -20.565 670.645 -20.235 ;
        RECT 668.955 -20.565 669.285 -20.235 ;
        RECT 667.595 -20.565 667.925 -20.235 ;
        RECT 666.235 -20.565 666.565 -20.235 ;
        RECT 664.875 -20.565 665.205 -20.235 ;
        RECT 663.515 -20.565 663.845 -20.235 ;
        RECT 659.435 -20.565 659.765 -20.235 ;
        RECT 656.715 -20.565 657.045 -20.235 ;
        RECT 655.355 -20.565 655.685 -20.235 ;
        RECT 653.995 -20.565 654.325 -20.235 ;
        RECT 652.635 -20.565 652.965 -20.235 ;
        RECT 651.275 -20.565 651.605 -20.235 ;
        RECT 649.915 -20.565 650.245 -20.235 ;
        RECT 648.555 -20.565 648.885 -20.235 ;
        RECT 643.115 -20.565 643.445 -20.235 ;
        RECT 641.755 -20.565 642.085 -20.235 ;
        RECT 640.395 -20.565 640.725 -20.235 ;
        RECT 639.035 -20.565 639.365 -20.235 ;
        RECT 637.675 -20.565 638.005 -20.235 ;
        RECT 636.315 -20.565 636.645 -20.235 ;
        RECT 634.955 -20.565 635.285 -20.235 ;
        RECT 633.595 -20.565 633.925 -20.235 ;
        RECT 628.155 -20.565 628.485 -20.235 ;
        RECT 626.795 -20.565 627.125 -20.235 ;
        RECT 625.435 -20.565 625.765 -20.235 ;
        RECT 624.075 -20.565 624.405 -20.235 ;
        RECT 622.715 -20.565 623.045 -20.235 ;
        RECT 621.355 -20.565 621.685 -20.235 ;
        RECT 619.995 -20.565 620.325 -20.235 ;
        RECT 618.635 -20.565 618.965 -20.235 ;
        RECT 613.195 -20.565 613.525 -20.235 ;
        RECT 611.835 -20.565 612.165 -20.235 ;
        RECT 610.475 -20.565 610.805 -20.235 ;
        RECT 609.115 -20.565 609.445 -20.235 ;
        RECT 607.755 -20.565 608.085 -20.235 ;
        RECT 606.395 -20.565 606.725 -20.235 ;
        RECT 605.035 -20.565 605.365 -20.235 ;
        RECT 603.675 -20.565 604.005 -20.235 ;
        RECT 598.235 -20.565 598.565 -20.235 ;
        RECT 596.875 -20.565 597.205 -20.235 ;
        RECT 595.515 -20.565 595.845 -20.235 ;
        RECT 594.155 -20.565 594.485 -20.235 ;
        RECT 592.795 -20.565 593.125 -20.235 ;
        RECT 591.435 -20.565 591.765 -20.235 ;
        RECT 590.075 -20.565 590.405 -20.235 ;
        RECT 588.715 -20.565 589.045 -20.235 ;
        RECT 583.275 -20.565 583.605 -20.235 ;
        RECT 581.915 -20.565 582.245 -20.235 ;
        RECT 580.555 -20.565 580.885 -20.235 ;
        RECT 579.195 -20.565 579.525 -20.235 ;
        RECT 577.835 -20.565 578.165 -20.235 ;
        RECT 576.475 -20.565 576.805 -20.235 ;
        RECT 575.115 -20.565 575.445 -20.235 ;
        RECT 573.755 -20.565 574.085 -20.235 ;
        RECT 568.315 -20.565 568.645 -20.235 ;
        RECT 566.955 -20.565 567.285 -20.235 ;
        RECT 565.595 -20.565 565.925 -20.235 ;
        RECT 564.235 -20.565 564.565 -20.235 ;
        RECT 562.875 -20.565 563.205 -20.235 ;
        RECT 561.515 -20.565 561.845 -20.235 ;
        RECT 560.155 -20.565 560.485 -20.235 ;
        RECT 558.795 -20.565 559.125 -20.235 ;
        RECT 553.355 -20.565 553.685 -20.235 ;
        RECT 551.995 -20.565 552.325 -20.235 ;
        RECT 550.635 -20.565 550.965 -20.235 ;
        RECT 549.275 -20.565 549.605 -20.235 ;
        RECT 547.915 -20.565 548.245 -20.235 ;
        RECT 546.555 -20.565 546.885 -20.235 ;
        RECT 545.195 -20.565 545.525 -20.235 ;
        RECT 543.835 -20.565 544.165 -20.235 ;
        RECT 538.395 -20.565 538.725 -20.235 ;
        RECT 537.035 -20.565 537.365 -20.235 ;
        RECT 535.675 -20.565 536.005 -20.235 ;
        RECT 534.315 -20.565 534.645 -20.235 ;
        RECT 532.955 -20.565 533.285 -20.235 ;
        RECT 531.595 -20.565 531.925 -20.235 ;
        RECT 530.235 -20.565 530.565 -20.235 ;
        RECT 528.875 -20.565 529.205 -20.235 ;
        RECT 523.435 -20.565 523.765 -20.235 ;
        RECT 522.075 -20.565 522.405 -20.235 ;
        RECT 520.715 -20.565 521.045 -20.235 ;
        RECT 519.355 -20.565 519.685 -20.235 ;
        RECT 517.995 -20.565 518.325 -20.235 ;
        RECT 516.635 -20.565 516.965 -20.235 ;
        RECT 515.275 -20.565 515.605 -20.235 ;
        RECT 513.915 -20.565 514.245 -20.235 ;
        RECT 508.475 -20.565 508.805 -20.235 ;
        RECT 507.115 -20.565 507.445 -20.235 ;
        RECT 505.755 -20.565 506.085 -20.235 ;
        RECT 504.395 -20.565 504.725 -20.235 ;
        RECT 503.035 -20.565 503.365 -20.235 ;
        RECT 501.675 -20.565 502.005 -20.235 ;
        RECT 500.315 -20.565 500.645 -20.235 ;
        RECT 498.955 -20.565 499.285 -20.235 ;
        RECT 493.515 -20.565 493.845 -20.235 ;
        RECT 492.155 -20.565 492.485 -20.235 ;
        RECT 490.795 -20.565 491.125 -20.235 ;
        RECT 489.435 -20.565 489.765 -20.235 ;
        RECT 488.075 -20.565 488.405 -20.235 ;
        RECT 486.715 -20.565 487.045 -20.235 ;
        RECT 485.355 -20.565 485.685 -20.235 ;
        RECT 483.995 -20.565 484.325 -20.235 ;
        RECT 478.555 -20.565 478.885 -20.235 ;
        RECT 477.195 -20.565 477.525 -20.235 ;
        RECT 475.835 -20.565 476.165 -20.235 ;
        RECT 474.475 -20.565 474.805 -20.235 ;
        RECT 473.115 -20.565 473.445 -20.235 ;
        RECT 471.755 -20.565 472.085 -20.235 ;
        RECT 470.395 -20.565 470.725 -20.235 ;
        RECT 469.035 -20.565 469.365 -20.235 ;
        RECT 463.595 -20.565 463.925 -20.235 ;
        RECT 462.235 -20.565 462.565 -20.235 ;
        RECT 460.875 -20.565 461.205 -20.235 ;
        RECT 459.515 -20.565 459.845 -20.235 ;
        RECT 458.155 -20.565 458.485 -20.235 ;
        RECT 456.795 -20.565 457.125 -20.235 ;
        RECT 455.435 -20.565 455.765 -20.235 ;
        RECT 454.075 -20.565 454.405 -20.235 ;
        RECT 448.635 -20.565 448.965 -20.235 ;
        RECT 447.275 -20.565 447.605 -20.235 ;
        RECT 445.915 -20.565 446.245 -20.235 ;
        RECT 444.555 -20.565 444.885 -20.235 ;
        RECT 443.195 -20.565 443.525 -20.235 ;
        RECT 441.835 -20.565 442.165 -20.235 ;
        RECT 440.475 -20.565 440.805 -20.235 ;
        RECT 439.115 -20.565 439.445 -20.235 ;
        RECT 436.395 -20.565 436.725 -20.235 ;
        RECT 433.675 -20.565 434.005 -20.235 ;
        RECT 432.315 -20.565 432.645 -20.235 ;
        RECT 430.955 -20.565 431.285 -20.235 ;
        RECT 429.595 -20.565 429.925 -20.235 ;
        RECT 428.235 -20.565 428.565 -20.235 ;
        RECT 426.875 -20.565 427.205 -20.235 ;
        RECT 425.515 -20.565 425.845 -20.235 ;
        RECT 424.155 -20.565 424.485 -20.235 ;
        RECT 421.435 -20.565 421.765 -20.235 ;
        RECT 418.715 -20.565 419.045 -20.235 ;
        RECT 417.355 -20.565 417.685 -20.235 ;
        RECT 415.995 -20.565 416.325 -20.235 ;
        RECT 414.635 -20.565 414.965 -20.235 ;
        RECT 413.275 -20.565 413.605 -20.235 ;
        RECT 411.915 -20.565 412.245 -20.235 ;
        RECT 410.555 -20.565 410.885 -20.235 ;
        RECT 406.475 -20.565 406.805 -20.235 ;
        RECT 403.755 -20.565 404.085 -20.235 ;
        RECT 402.395 -20.565 402.725 -20.235 ;
        RECT 401.035 -20.565 401.365 -20.235 ;
        RECT 399.675 -20.565 400.005 -20.235 ;
        RECT 398.315 -20.565 398.645 -20.235 ;
        RECT 396.955 -20.565 397.285 -20.235 ;
        RECT 395.595 -20.565 395.925 -20.235 ;
        RECT 391.515 -20.565 391.845 -20.235 ;
        RECT 388.795 -20.565 389.125 -20.235 ;
        RECT 387.435 -20.565 387.765 -20.235 ;
        RECT 386.075 -20.565 386.405 -20.235 ;
        RECT 384.715 -20.565 385.045 -20.235 ;
        RECT 383.355 -20.565 383.685 -20.235 ;
        RECT 381.995 -20.565 382.325 -20.235 ;
        RECT 380.635 -20.565 380.965 -20.235 ;
        RECT 376.555 -20.565 376.885 -20.235 ;
        RECT 373.835 -20.565 374.165 -20.235 ;
        RECT 372.475 -20.565 372.805 -20.235 ;
        RECT 371.115 -20.565 371.445 -20.235 ;
        RECT 369.755 -20.565 370.085 -20.235 ;
        RECT 368.395 -20.565 368.725 -20.235 ;
        RECT 367.035 -20.565 367.365 -20.235 ;
        RECT 365.675 -20.565 366.005 -20.235 ;
        RECT 361.595 -20.565 361.925 -20.235 ;
        RECT 358.875 -20.565 359.205 -20.235 ;
        RECT 357.515 -20.565 357.845 -20.235 ;
        RECT 356.155 -20.565 356.485 -20.235 ;
        RECT 354.795 -20.565 355.125 -20.235 ;
        RECT 353.435 -20.565 353.765 -20.235 ;
        RECT 352.075 -20.565 352.405 -20.235 ;
        RECT 350.715 -20.565 351.045 -20.235 ;
        RECT 346.635 -20.565 346.965 -20.235 ;
        RECT 343.915 -20.565 344.245 -20.235 ;
        RECT 342.555 -20.565 342.885 -20.235 ;
        RECT 341.195 -20.565 341.525 -20.235 ;
        RECT 339.835 -20.565 340.165 -20.235 ;
        RECT 338.475 -20.565 338.805 -20.235 ;
        RECT 337.115 -20.565 337.445 -20.235 ;
        RECT 335.755 -20.565 336.085 -20.235 ;
        RECT 331.675 -20.565 332.005 -20.235 ;
        RECT 328.955 -20.565 329.285 -20.235 ;
        RECT 327.595 -20.565 327.925 -20.235 ;
        RECT 326.235 -20.565 326.565 -20.235 ;
        RECT 324.875 -20.565 325.205 -20.235 ;
        RECT 323.515 -20.565 323.845 -20.235 ;
        RECT 322.155 -20.565 322.485 -20.235 ;
        RECT 320.795 -20.565 321.125 -20.235 ;
        RECT 316.715 -20.565 317.045 -20.235 ;
        RECT 313.995 -20.565 314.325 -20.235 ;
        RECT 312.635 -20.565 312.965 -20.235 ;
        RECT 311.275 -20.565 311.605 -20.235 ;
        RECT 309.915 -20.565 310.245 -20.235 ;
        RECT 308.555 -20.565 308.885 -20.235 ;
        RECT 307.195 -20.565 307.525 -20.235 ;
        RECT 305.835 -20.565 306.165 -20.235 ;
        RECT 300.395 -20.565 300.725 -20.235 ;
        RECT 299.035 -20.565 299.365 -20.235 ;
        RECT 297.675 -20.565 298.005 -20.235 ;
        RECT 296.315 -20.565 296.645 -20.235 ;
        RECT 294.955 -20.565 295.285 -20.235 ;
        RECT 293.595 -20.565 293.925 -20.235 ;
        RECT 292.235 -20.565 292.565 -20.235 ;
        RECT 290.875 -20.565 291.205 -20.235 ;
        RECT 285.435 -20.565 285.765 -20.235 ;
        RECT 284.075 -20.565 284.405 -20.235 ;
        RECT 282.715 -20.565 283.045 -20.235 ;
        RECT 281.355 -20.565 281.685 -20.235 ;
        RECT 279.995 -20.565 280.325 -20.235 ;
        RECT 278.635 -20.565 278.965 -20.235 ;
        RECT 277.275 -20.565 277.605 -20.235 ;
        RECT 275.915 -20.565 276.245 -20.235 ;
        RECT 270.475 -20.565 270.805 -20.235 ;
        RECT 269.115 -20.565 269.445 -20.235 ;
        RECT 267.755 -20.565 268.085 -20.235 ;
        RECT 266.395 -20.565 266.725 -20.235 ;
        RECT 265.035 -20.565 265.365 -20.235 ;
        RECT 263.675 -20.565 264.005 -20.235 ;
        RECT 262.315 -20.565 262.645 -20.235 ;
        RECT 260.955 -20.565 261.285 -20.235 ;
        RECT 255.515 -20.565 255.845 -20.235 ;
        RECT 254.155 -20.565 254.485 -20.235 ;
        RECT 252.795 -20.565 253.125 -20.235 ;
        RECT 251.435 -20.565 251.765 -20.235 ;
        RECT 250.075 -20.565 250.405 -20.235 ;
        RECT 248.715 -20.565 249.045 -20.235 ;
        RECT 247.355 -20.565 247.685 -20.235 ;
        RECT 245.995 -20.565 246.325 -20.235 ;
        RECT 240.555 -20.565 240.885 -20.235 ;
        RECT 239.195 -20.565 239.525 -20.235 ;
        RECT 237.835 -20.565 238.165 -20.235 ;
        RECT 236.475 -20.565 236.805 -20.235 ;
        RECT 235.115 -20.565 235.445 -20.235 ;
        RECT 233.755 -20.565 234.085 -20.235 ;
        RECT 232.395 -20.565 232.725 -20.235 ;
        RECT 231.035 -20.565 231.365 -20.235 ;
        RECT 225.595 -20.565 225.925 -20.235 ;
        RECT 224.235 -20.565 224.565 -20.235 ;
        RECT 222.875 -20.565 223.205 -20.235 ;
        RECT 221.515 -20.565 221.845 -20.235 ;
        RECT 220.155 -20.565 220.485 -20.235 ;
        RECT 218.795 -20.565 219.125 -20.235 ;
        RECT 217.435 -20.565 217.765 -20.235 ;
        RECT 216.075 -20.565 216.405 -20.235 ;
        RECT 210.635 -20.565 210.965 -20.235 ;
        RECT 209.275 -20.565 209.605 -20.235 ;
        RECT 207.915 -20.565 208.245 -20.235 ;
        RECT 206.555 -20.565 206.885 -20.235 ;
        RECT 205.195 -20.565 205.525 -20.235 ;
        RECT 203.835 -20.565 204.165 -20.235 ;
        RECT 202.475 -20.565 202.805 -20.235 ;
        RECT 201.115 -20.565 201.445 -20.235 ;
        RECT 195.675 -20.565 196.005 -20.235 ;
        RECT 194.315 -20.565 194.645 -20.235 ;
        RECT 192.955 -20.565 193.285 -20.235 ;
        RECT 191.595 -20.565 191.925 -20.235 ;
        RECT 190.235 -20.565 190.565 -20.235 ;
        RECT 188.875 -20.565 189.205 -20.235 ;
        RECT 187.515 -20.565 187.845 -20.235 ;
        RECT 186.155 -20.565 186.485 -20.235 ;
        RECT 180.715 -20.565 181.045 -20.235 ;
        RECT 179.355 -20.565 179.685 -20.235 ;
        RECT 177.995 -20.565 178.325 -20.235 ;
        RECT 176.635 -20.565 176.965 -20.235 ;
        RECT 175.275 -20.565 175.605 -20.235 ;
        RECT 173.915 -20.565 174.245 -20.235 ;
        RECT 172.555 -20.565 172.885 -20.235 ;
        RECT 171.195 -20.565 171.525 -20.235 ;
        RECT 165.755 -20.565 166.085 -20.235 ;
        RECT 164.395 -20.565 164.725 -20.235 ;
        RECT 163.035 -20.565 163.365 -20.235 ;
        RECT 161.675 -20.565 162.005 -20.235 ;
        RECT 160.315 -20.565 160.645 -20.235 ;
        RECT 158.955 -20.565 159.285 -20.235 ;
        RECT 157.595 -20.565 157.925 -20.235 ;
        RECT 156.235 -20.565 156.565 -20.235 ;
        RECT 150.795 -20.565 151.125 -20.235 ;
        RECT 149.435 -20.565 149.765 -20.235 ;
        RECT 148.075 -20.565 148.405 -20.235 ;
        RECT 146.715 -20.565 147.045 -20.235 ;
        RECT 145.355 -20.565 145.685 -20.235 ;
        RECT 143.995 -20.565 144.325 -20.235 ;
        RECT 142.635 -20.565 142.965 -20.235 ;
        RECT 141.275 -20.565 141.605 -20.235 ;
        RECT 135.835 -20.565 136.165 -20.235 ;
        RECT 134.475 -20.565 134.805 -20.235 ;
        RECT 133.115 -20.565 133.445 -20.235 ;
        RECT 131.755 -20.565 132.085 -20.235 ;
        RECT 130.395 -20.565 130.725 -20.235 ;
        RECT 129.035 -20.565 129.365 -20.235 ;
        RECT 127.675 -20.565 128.005 -20.235 ;
        RECT 126.315 -20.565 126.645 -20.235 ;
        RECT 120.875 -20.565 121.205 -20.235 ;
        RECT 119.515 -20.565 119.845 -20.235 ;
        RECT 118.155 -20.565 118.485 -20.235 ;
        RECT 116.795 -20.565 117.125 -20.235 ;
        RECT 115.435 -20.565 115.765 -20.235 ;
        RECT 114.075 -20.565 114.405 -20.235 ;
        RECT 112.715 -20.565 113.045 -20.235 ;
        RECT 111.355 -20.565 111.685 -20.235 ;
        RECT 105.915 -20.565 106.245 -20.235 ;
        RECT 104.555 -20.565 104.885 -20.235 ;
        RECT 103.195 -20.565 103.525 -20.235 ;
        RECT 101.835 -20.565 102.165 -20.235 ;
        RECT 100.475 -20.565 100.805 -20.235 ;
        RECT 99.115 -20.565 99.445 -20.235 ;
        RECT 97.755 -20.565 98.085 -20.235 ;
        RECT 96.395 -20.565 96.725 -20.235 ;
        RECT 93.675 -20.565 94.005 -20.235 ;
        RECT 90.955 -20.565 91.285 -20.235 ;
        RECT 89.595 -20.565 89.925 -20.235 ;
        RECT 88.235 -20.565 88.565 -20.235 ;
        RECT 86.875 -20.565 87.205 -20.235 ;
        RECT 85.515 -20.565 85.845 -20.235 ;
        RECT 84.155 -20.565 84.485 -20.235 ;
        RECT 82.795 -20.565 83.125 -20.235 ;
        RECT 81.435 -20.565 81.765 -20.235 ;
        RECT 78.715 -20.565 79.045 -20.235 ;
        RECT 75.995 -20.565 76.325 -20.235 ;
        RECT 74.635 -20.565 74.965 -20.235 ;
        RECT 73.275 -20.565 73.605 -20.235 ;
        RECT 71.915 -20.565 72.245 -20.235 ;
        RECT 70.555 -20.565 70.885 -20.235 ;
        RECT 69.195 -20.565 69.525 -20.235 ;
        RECT 67.835 -20.565 68.165 -20.235 ;
        RECT 63.755 -20.565 64.085 -20.235 ;
        RECT 61.035 -20.565 61.365 -20.235 ;
        RECT 59.675 -20.565 60.005 -20.235 ;
        RECT 58.315 -20.565 58.645 -20.235 ;
        RECT 56.955 -20.565 57.285 -20.235 ;
        RECT 55.595 -20.565 55.925 -20.235 ;
        RECT 54.235 -20.565 54.565 -20.235 ;
        RECT 52.875 -20.565 53.205 -20.235 ;
        RECT 48.795 -20.565 49.125 -20.235 ;
        RECT 46.075 -20.565 46.405 -20.235 ;
        RECT 44.715 -20.565 45.045 -20.235 ;
        RECT 43.355 -20.565 43.685 -20.235 ;
        RECT 41.995 -20.565 42.325 -20.235 ;
        RECT 40.635 -20.565 40.965 -20.235 ;
        RECT 39.275 -20.565 39.605 -20.235 ;
        RECT 37.915 -20.565 38.245 -20.235 ;
        RECT 33.835 -20.565 34.165 -20.235 ;
        RECT 31.115 -20.565 31.445 -20.235 ;
        RECT 29.755 -20.565 30.085 -20.235 ;
        RECT 28.395 -20.565 28.725 -20.235 ;
        RECT 27.035 -20.565 27.365 -20.235 ;
        RECT 25.675 -20.565 26.005 -20.235 ;
        RECT 24.315 -20.565 24.645 -20.235 ;
        RECT 22.955 -20.565 23.285 -20.235 ;
        RECT 18.875 -20.565 19.205 -20.235 ;
        RECT 16.155 -20.565 16.485 -20.235 ;
        RECT 14.795 -20.565 15.125 -20.235 ;
        RECT 13.435 -20.565 13.765 -20.235 ;
        RECT 12.075 -20.565 12.405 -20.235 ;
        RECT 10.715 -20.565 11.045 -20.235 ;
        RECT 9.355 -20.565 9.685 -20.235 ;
        RECT 7.995 -20.565 8.325 -20.235 ;
        RECT 6.635 -20.565 6.965 -20.235 ;
        RECT 3.915 -20.565 4.245 -20.235 ;
        RECT 2.555 -20.565 2.885 -20.235 ;
        RECT 1.195 -20.565 1.525 -20.235 ;
        RECT -0.165 -20.565 0.165 -20.235 ;
        RECT -1.525 -20.565 -1.195 -20.235 ;
        RECT 954.555 -20.565 954.885 -20.235 ;
        RECT 920.555 -20.56 954.885 -20.24 ;
        RECT 953.195 -20.565 953.525 -20.235 ;
        RECT 951.835 -20.565 952.165 -20.235 ;
        RECT 950.475 -20.565 950.805 -20.235 ;
        RECT 949.115 -20.565 949.445 -20.235 ;
        RECT 947.755 -20.565 948.085 -20.235 ;
        RECT 946.395 -20.565 946.725 -20.235 ;
        RECT 945.035 -20.565 945.365 -20.235 ;
        RECT 940.955 -20.565 941.285 -20.235 ;
        RECT 939.595 -20.565 939.925 -20.235 ;
        RECT 938.235 -20.565 938.565 -20.235 ;
        RECT 936.875 -20.565 937.205 -20.235 ;
        RECT 935.515 -20.565 935.845 -20.235 ;
        RECT 934.155 -20.565 934.485 -20.235 ;
        RECT 932.795 -20.565 933.125 -20.235 ;
        RECT 931.435 -20.565 931.765 -20.235 ;
        RECT 925.995 -20.565 926.325 -20.235 ;
        RECT 924.635 -20.565 924.965 -20.235 ;
        RECT 923.275 -20.565 923.605 -20.235 ;
        RECT 921.915 -20.565 922.245 -20.235 ;
        RECT 920.555 -20.565 920.885 -20.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 919.88 -30.08 926.32 -29.76 ;
        RECT 924.635 -30.085 924.965 -29.755 ;
        RECT 923.275 -30.085 923.605 -29.755 ;
        RECT 921.915 -30.085 922.245 -29.755 ;
        RECT 920.555 -30.085 920.885 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 920.555 -23.285 920.885 -22.955 ;
        RECT 916.475 -23.285 916.805 -22.955 ;
        RECT 915.8 -23.28 927 -22.96 ;
        RECT 924.635 -23.285 924.965 -22.955 ;
        RECT 923.275 -23.285 923.605 -22.955 ;
        RECT 921.915 -23.285 922.245 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.88 -30.08 687.64 -29.76 ;
        RECT 686.635 -30.085 686.965 -29.755 ;
        RECT 685.275 -30.085 685.605 -29.755 ;
        RECT 683.915 -30.085 684.245 -29.755 ;
        RECT 682.555 -30.085 682.885 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.12 -23.28 688.32 -22.96 ;
        RECT 686.635 -23.285 686.965 -22.955 ;
        RECT 685.275 -23.285 685.605 -22.955 ;
        RECT 683.915 -23.285 684.245 -22.955 ;
        RECT 682.555 -23.285 682.885 -22.955 ;
        RECT 678.475 -23.285 678.805 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 677.8 -27.36 688.32 -27.04 ;
        RECT 686.635 -27.365 686.965 -27.035 ;
        RECT 685.275 -27.365 685.605 -27.035 ;
        RECT 683.915 -27.365 684.245 -27.035 ;
        RECT 682.555 -27.365 682.885 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 687.995 -35.525 688.325 -35.195 ;
        RECT 681.88 -35.52 688.325 -35.2 ;
        RECT 686.635 -35.525 686.965 -35.195 ;
        RECT 685.275 -35.525 685.605 -35.195 ;
        RECT 683.915 -35.525 684.245 -35.195 ;
        RECT 682.555 -35.525 682.885 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 681.88 -26 692.4 -25.68 ;
        RECT 690.715 -26.005 691.045 -25.675 ;
        RECT 689.355 -26.005 689.685 -25.675 ;
        RECT 686.635 -26.005 686.965 -25.675 ;
        RECT 685.275 -26.005 685.605 -25.675 ;
        RECT 683.915 -26.005 684.245 -25.675 ;
        RECT 682.555 -26.005 682.885 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.16 -30.08 702.6 -29.76 ;
        RECT 701.595 -30.085 701.925 -29.755 ;
        RECT 700.235 -30.085 700.565 -29.755 ;
        RECT 698.875 -30.085 699.205 -29.755 ;
        RECT 697.515 -30.085 697.845 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.08 -23.28 703.28 -22.96 ;
        RECT 701.595 -23.285 701.925 -22.955 ;
        RECT 700.235 -23.285 700.565 -22.955 ;
        RECT 698.875 -23.285 699.205 -22.955 ;
        RECT 697.515 -23.285 697.845 -22.955 ;
        RECT 696.155 -23.285 696.485 -22.955 ;
        RECT 693.435 -23.285 693.765 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 692.76 -27.36 703.28 -27.04 ;
        RECT 701.595 -27.365 701.925 -27.035 ;
        RECT 700.235 -27.365 700.565 -27.035 ;
        RECT 698.875 -27.365 699.205 -27.035 ;
        RECT 697.515 -27.365 697.845 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 702.955 -35.525 703.285 -35.195 ;
        RECT 696.16 -35.52 703.285 -35.2 ;
        RECT 701.595 -35.525 701.925 -35.195 ;
        RECT 700.235 -35.525 700.565 -35.195 ;
        RECT 698.875 -35.525 699.205 -35.195 ;
        RECT 697.515 -35.525 697.845 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 696.16 -26 707.36 -25.68 ;
        RECT 705.675 -26.005 706.005 -25.675 ;
        RECT 704.315 -26.005 704.645 -25.675 ;
        RECT 701.595 -26.005 701.925 -25.675 ;
        RECT 700.235 -26.005 700.565 -25.675 ;
        RECT 698.875 -26.005 699.205 -25.675 ;
        RECT 697.515 -26.005 697.845 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.12 -30.08 717.56 -29.76 ;
        RECT 716.555 -30.085 716.885 -29.755 ;
        RECT 715.195 -30.085 715.525 -29.755 ;
        RECT 713.835 -30.085 714.165 -29.755 ;
        RECT 712.475 -30.085 712.805 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.04 -23.28 718.24 -22.96 ;
        RECT 716.555 -23.285 716.885 -22.955 ;
        RECT 715.195 -23.285 715.525 -22.955 ;
        RECT 713.835 -23.285 714.165 -22.955 ;
        RECT 712.475 -23.285 712.805 -22.955 ;
        RECT 711.115 -23.285 711.445 -22.955 ;
        RECT 708.395 -23.285 708.725 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 707.72 -27.36 718.24 -27.04 ;
        RECT 716.555 -27.365 716.885 -27.035 ;
        RECT 715.195 -27.365 715.525 -27.035 ;
        RECT 713.835 -27.365 714.165 -27.035 ;
        RECT 712.475 -27.365 712.805 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 717.915 -35.525 718.245 -35.195 ;
        RECT 711.12 -35.52 718.245 -35.2 ;
        RECT 716.555 -35.525 716.885 -35.195 ;
        RECT 715.195 -35.525 715.525 -35.195 ;
        RECT 713.835 -35.525 714.165 -35.195 ;
        RECT 712.475 -35.525 712.805 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 711.12 -26 722.32 -25.68 ;
        RECT 720.635 -26.005 720.965 -25.675 ;
        RECT 719.275 -26.005 719.605 -25.675 ;
        RECT 716.555 -26.005 716.885 -25.675 ;
        RECT 715.195 -26.005 715.525 -25.675 ;
        RECT 713.835 -26.005 714.165 -25.675 ;
        RECT 712.475 -26.005 712.805 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.08 -30.08 732.52 -29.76 ;
        RECT 731.515 -30.085 731.845 -29.755 ;
        RECT 730.155 -30.085 730.485 -29.755 ;
        RECT 728.795 -30.085 729.125 -29.755 ;
        RECT 727.435 -30.085 727.765 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 722 -23.28 733.2 -22.96 ;
        RECT 731.515 -23.285 731.845 -22.955 ;
        RECT 730.155 -23.285 730.485 -22.955 ;
        RECT 728.795 -23.285 729.125 -22.955 ;
        RECT 727.435 -23.285 727.765 -22.955 ;
        RECT 726.075 -23.285 726.405 -22.955 ;
        RECT 723.355 -23.285 723.685 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 722.68 -27.36 733.2 -27.04 ;
        RECT 731.515 -27.365 731.845 -27.035 ;
        RECT 730.155 -27.365 730.485 -27.035 ;
        RECT 728.795 -27.365 729.125 -27.035 ;
        RECT 727.435 -27.365 727.765 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 732.875 -35.525 733.205 -35.195 ;
        RECT 726.08 -35.52 733.205 -35.2 ;
        RECT 731.515 -35.525 731.845 -35.195 ;
        RECT 730.155 -35.525 730.485 -35.195 ;
        RECT 728.795 -35.525 729.125 -35.195 ;
        RECT 727.435 -35.525 727.765 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 726.08 -26 736.6 -25.68 ;
        RECT 735.595 -26.005 735.925 -25.675 ;
        RECT 734.235 -26.005 734.565 -25.675 ;
        RECT 731.515 -26.005 731.845 -25.675 ;
        RECT 730.155 -26.005 730.485 -25.675 ;
        RECT 728.795 -26.005 729.125 -25.675 ;
        RECT 727.435 -26.005 727.765 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -17.84 743.755 -17.52 ;
        RECT 742.395 -17.845 742.725 -17.515 ;
        RECT 741.035 -17.845 741.365 -17.515 ;
        RECT 739.675 -17.845 740.005 -17.515 ;
        RECT 738.315 -17.845 738.645 -17.515 ;
        RECT 735.595 -17.845 735.925 -17.515 ;
        RECT 734.235 -17.845 734.565 -17.515 ;
        RECT 732.875 -17.845 733.205 -17.515 ;
        RECT 731.515 -17.845 731.845 -17.515 ;
        RECT 730.155 -17.845 730.485 -17.515 ;
        RECT 728.795 -17.845 729.125 -17.515 ;
        RECT 727.435 -17.845 727.765 -17.515 ;
        RECT 726.075 -17.845 726.405 -17.515 ;
        RECT 724.715 -17.845 725.045 -17.515 ;
        RECT 723.355 -17.845 723.685 -17.515 ;
        RECT 720.635 -17.845 720.965 -17.515 ;
        RECT 719.275 -17.845 719.605 -17.515 ;
        RECT 717.915 -17.845 718.245 -17.515 ;
        RECT 716.555 -17.845 716.885 -17.515 ;
        RECT 715.195 -17.845 715.525 -17.515 ;
        RECT 713.835 -17.845 714.165 -17.515 ;
        RECT 712.475 -17.845 712.805 -17.515 ;
        RECT 711.115 -17.845 711.445 -17.515 ;
        RECT 709.755 -17.845 710.085 -17.515 ;
        RECT 708.395 -17.845 708.725 -17.515 ;
        RECT 705.675 -17.845 706.005 -17.515 ;
        RECT 704.315 -17.845 704.645 -17.515 ;
        RECT 702.955 -17.845 703.285 -17.515 ;
        RECT 701.595 -17.845 701.925 -17.515 ;
        RECT 700.235 -17.845 700.565 -17.515 ;
        RECT 698.875 -17.845 699.205 -17.515 ;
        RECT 697.515 -17.845 697.845 -17.515 ;
        RECT 696.155 -17.845 696.485 -17.515 ;
        RECT 694.795 -17.845 695.125 -17.515 ;
        RECT 693.435 -17.845 693.765 -17.515 ;
        RECT 690.715 -17.845 691.045 -17.515 ;
        RECT 689.355 -17.845 689.685 -17.515 ;
        RECT 687.995 -17.845 688.325 -17.515 ;
        RECT 686.635 -17.845 686.965 -17.515 ;
        RECT 685.275 -17.845 685.605 -17.515 ;
        RECT 683.915 -17.845 684.245 -17.515 ;
        RECT 682.555 -17.845 682.885 -17.515 ;
        RECT 681.195 -17.845 681.525 -17.515 ;
        RECT 679.835 -17.845 680.165 -17.515 ;
        RECT 678.475 -17.845 678.805 -17.515 ;
        RECT 675.755 -17.845 676.085 -17.515 ;
        RECT 674.395 -17.845 674.725 -17.515 ;
        RECT 673.035 -17.845 673.365 -17.515 ;
        RECT 671.675 -17.845 672.005 -17.515 ;
        RECT 670.315 -17.845 670.645 -17.515 ;
        RECT 668.955 -17.845 669.285 -17.515 ;
        RECT 667.595 -17.845 667.925 -17.515 ;
        RECT 666.235 -17.845 666.565 -17.515 ;
        RECT 664.875 -17.845 665.205 -17.515 ;
        RECT 663.515 -17.845 663.845 -17.515 ;
        RECT 660.795 -17.845 661.125 -17.515 ;
        RECT 659.435 -17.845 659.765 -17.515 ;
        RECT 658.075 -17.845 658.405 -17.515 ;
        RECT 656.715 -17.845 657.045 -17.515 ;
        RECT 655.355 -17.845 655.685 -17.515 ;
        RECT 653.995 -17.845 654.325 -17.515 ;
        RECT 652.635 -17.845 652.965 -17.515 ;
        RECT 651.275 -17.845 651.605 -17.515 ;
        RECT 649.915 -17.845 650.245 -17.515 ;
        RECT 648.555 -17.845 648.885 -17.515 ;
        RECT 645.835 -17.845 646.165 -17.515 ;
        RECT 644.475 -17.845 644.805 -17.515 ;
        RECT 643.115 -17.845 643.445 -17.515 ;
        RECT 641.755 -17.845 642.085 -17.515 ;
        RECT 640.395 -17.845 640.725 -17.515 ;
        RECT 639.035 -17.845 639.365 -17.515 ;
        RECT 637.675 -17.845 638.005 -17.515 ;
        RECT 636.315 -17.845 636.645 -17.515 ;
        RECT 634.955 -17.845 635.285 -17.515 ;
        RECT 633.595 -17.845 633.925 -17.515 ;
        RECT 630.875 -17.845 631.205 -17.515 ;
        RECT 629.515 -17.845 629.845 -17.515 ;
        RECT 628.155 -17.845 628.485 -17.515 ;
        RECT 626.795 -17.845 627.125 -17.515 ;
        RECT 625.435 -17.845 625.765 -17.515 ;
        RECT 624.075 -17.845 624.405 -17.515 ;
        RECT 622.715 -17.845 623.045 -17.515 ;
        RECT 621.355 -17.845 621.685 -17.515 ;
        RECT 619.995 -17.845 620.325 -17.515 ;
        RECT 618.635 -17.845 618.965 -17.515 ;
        RECT 615.915 -17.845 616.245 -17.515 ;
        RECT 614.555 -17.845 614.885 -17.515 ;
        RECT 613.195 -17.845 613.525 -17.515 ;
        RECT 611.835 -17.845 612.165 -17.515 ;
        RECT 610.475 -17.845 610.805 -17.515 ;
        RECT 609.115 -17.845 609.445 -17.515 ;
        RECT 607.755 -17.845 608.085 -17.515 ;
        RECT 606.395 -17.845 606.725 -17.515 ;
        RECT 605.035 -17.845 605.365 -17.515 ;
        RECT 603.675 -17.845 604.005 -17.515 ;
        RECT 600.955 -17.845 601.285 -17.515 ;
        RECT 599.595 -17.845 599.925 -17.515 ;
        RECT 598.235 -17.845 598.565 -17.515 ;
        RECT 596.875 -17.845 597.205 -17.515 ;
        RECT 595.515 -17.845 595.845 -17.515 ;
        RECT 594.155 -17.845 594.485 -17.515 ;
        RECT 592.795 -17.845 593.125 -17.515 ;
        RECT 591.435 -17.845 591.765 -17.515 ;
        RECT 590.075 -17.845 590.405 -17.515 ;
        RECT 588.715 -17.845 589.045 -17.515 ;
        RECT 585.995 -17.845 586.325 -17.515 ;
        RECT 584.635 -17.845 584.965 -17.515 ;
        RECT 583.275 -17.845 583.605 -17.515 ;
        RECT 581.915 -17.845 582.245 -17.515 ;
        RECT 580.555 -17.845 580.885 -17.515 ;
        RECT 579.195 -17.845 579.525 -17.515 ;
        RECT 577.835 -17.845 578.165 -17.515 ;
        RECT 576.475 -17.845 576.805 -17.515 ;
        RECT 575.115 -17.845 575.445 -17.515 ;
        RECT 573.755 -17.845 574.085 -17.515 ;
        RECT 571.035 -17.845 571.365 -17.515 ;
        RECT 569.675 -17.845 570.005 -17.515 ;
        RECT 568.315 -17.845 568.645 -17.515 ;
        RECT 566.955 -17.845 567.285 -17.515 ;
        RECT 565.595 -17.845 565.925 -17.515 ;
        RECT 564.235 -17.845 564.565 -17.515 ;
        RECT 562.875 -17.845 563.205 -17.515 ;
        RECT 561.515 -17.845 561.845 -17.515 ;
        RECT 560.155 -17.845 560.485 -17.515 ;
        RECT 558.795 -17.845 559.125 -17.515 ;
        RECT 556.075 -17.845 556.405 -17.515 ;
        RECT 554.715 -17.845 555.045 -17.515 ;
        RECT 553.355 -17.845 553.685 -17.515 ;
        RECT 551.995 -17.845 552.325 -17.515 ;
        RECT 550.635 -17.845 550.965 -17.515 ;
        RECT 549.275 -17.845 549.605 -17.515 ;
        RECT 547.915 -17.845 548.245 -17.515 ;
        RECT 546.555 -17.845 546.885 -17.515 ;
        RECT 545.195 -17.845 545.525 -17.515 ;
        RECT 543.835 -17.845 544.165 -17.515 ;
        RECT 541.115 -17.845 541.445 -17.515 ;
        RECT 539.755 -17.845 540.085 -17.515 ;
        RECT 538.395 -17.845 538.725 -17.515 ;
        RECT 537.035 -17.845 537.365 -17.515 ;
        RECT 535.675 -17.845 536.005 -17.515 ;
        RECT 534.315 -17.845 534.645 -17.515 ;
        RECT 532.955 -17.845 533.285 -17.515 ;
        RECT 531.595 -17.845 531.925 -17.515 ;
        RECT 530.235 -17.845 530.565 -17.515 ;
        RECT 528.875 -17.845 529.205 -17.515 ;
        RECT 526.155 -17.845 526.485 -17.515 ;
        RECT 524.795 -17.845 525.125 -17.515 ;
        RECT 523.435 -17.845 523.765 -17.515 ;
        RECT 522.075 -17.845 522.405 -17.515 ;
        RECT 520.715 -17.845 521.045 -17.515 ;
        RECT 519.355 -17.845 519.685 -17.515 ;
        RECT 517.995 -17.845 518.325 -17.515 ;
        RECT 516.635 -17.845 516.965 -17.515 ;
        RECT 515.275 -17.845 515.605 -17.515 ;
        RECT 513.915 -17.845 514.245 -17.515 ;
        RECT 511.195 -17.845 511.525 -17.515 ;
        RECT 509.835 -17.845 510.165 -17.515 ;
        RECT 508.475 -17.845 508.805 -17.515 ;
        RECT 507.115 -17.845 507.445 -17.515 ;
        RECT 505.755 -17.845 506.085 -17.515 ;
        RECT 504.395 -17.845 504.725 -17.515 ;
        RECT 503.035 -17.845 503.365 -17.515 ;
        RECT 501.675 -17.845 502.005 -17.515 ;
        RECT 500.315 -17.845 500.645 -17.515 ;
        RECT 498.955 -17.845 499.285 -17.515 ;
        RECT 496.235 -17.845 496.565 -17.515 ;
        RECT 494.875 -17.845 495.205 -17.515 ;
        RECT 493.515 -17.845 493.845 -17.515 ;
        RECT 492.155 -17.845 492.485 -17.515 ;
        RECT 490.795 -17.845 491.125 -17.515 ;
        RECT 489.435 -17.845 489.765 -17.515 ;
        RECT 488.075 -17.845 488.405 -17.515 ;
        RECT 486.715 -17.845 487.045 -17.515 ;
        RECT 485.355 -17.845 485.685 -17.515 ;
        RECT 483.995 -17.845 484.325 -17.515 ;
        RECT 481.275 -17.845 481.605 -17.515 ;
        RECT 479.915 -17.845 480.245 -17.515 ;
        RECT 478.555 -17.845 478.885 -17.515 ;
        RECT 477.195 -17.845 477.525 -17.515 ;
        RECT 475.835 -17.845 476.165 -17.515 ;
        RECT 474.475 -17.845 474.805 -17.515 ;
        RECT 473.115 -17.845 473.445 -17.515 ;
        RECT 471.755 -17.845 472.085 -17.515 ;
        RECT 470.395 -17.845 470.725 -17.515 ;
        RECT 469.035 -17.845 469.365 -17.515 ;
        RECT 466.315 -17.845 466.645 -17.515 ;
        RECT 464.955 -17.845 465.285 -17.515 ;
        RECT 463.595 -17.845 463.925 -17.515 ;
        RECT 462.235 -17.845 462.565 -17.515 ;
        RECT 460.875 -17.845 461.205 -17.515 ;
        RECT 459.515 -17.845 459.845 -17.515 ;
        RECT 458.155 -17.845 458.485 -17.515 ;
        RECT 456.795 -17.845 457.125 -17.515 ;
        RECT 455.435 -17.845 455.765 -17.515 ;
        RECT 454.075 -17.845 454.405 -17.515 ;
        RECT 451.355 -17.845 451.685 -17.515 ;
        RECT 449.995 -17.845 450.325 -17.515 ;
        RECT 448.635 -17.845 448.965 -17.515 ;
        RECT 447.275 -17.845 447.605 -17.515 ;
        RECT 445.915 -17.845 446.245 -17.515 ;
        RECT 444.555 -17.845 444.885 -17.515 ;
        RECT 443.195 -17.845 443.525 -17.515 ;
        RECT 441.835 -17.845 442.165 -17.515 ;
        RECT 440.475 -17.845 440.805 -17.515 ;
        RECT 439.115 -17.845 439.445 -17.515 ;
        RECT 436.395 -17.845 436.725 -17.515 ;
        RECT 435.035 -17.845 435.365 -17.515 ;
        RECT 433.675 -17.845 434.005 -17.515 ;
        RECT 432.315 -17.845 432.645 -17.515 ;
        RECT 430.955 -17.845 431.285 -17.515 ;
        RECT 429.595 -17.845 429.925 -17.515 ;
        RECT 428.235 -17.845 428.565 -17.515 ;
        RECT 426.875 -17.845 427.205 -17.515 ;
        RECT 425.515 -17.845 425.845 -17.515 ;
        RECT 424.155 -17.845 424.485 -17.515 ;
        RECT 421.435 -17.845 421.765 -17.515 ;
        RECT 420.075 -17.845 420.405 -17.515 ;
        RECT 418.715 -17.845 419.045 -17.515 ;
        RECT 417.355 -17.845 417.685 -17.515 ;
        RECT 415.995 -17.845 416.325 -17.515 ;
        RECT 414.635 -17.845 414.965 -17.515 ;
        RECT 413.275 -17.845 413.605 -17.515 ;
        RECT 411.915 -17.845 412.245 -17.515 ;
        RECT 410.555 -17.845 410.885 -17.515 ;
        RECT 407.835 -17.845 408.165 -17.515 ;
        RECT 406.475 -17.845 406.805 -17.515 ;
        RECT 405.115 -17.845 405.445 -17.515 ;
        RECT 403.755 -17.845 404.085 -17.515 ;
        RECT 402.395 -17.845 402.725 -17.515 ;
        RECT 401.035 -17.845 401.365 -17.515 ;
        RECT 399.675 -17.845 400.005 -17.515 ;
        RECT 398.315 -17.845 398.645 -17.515 ;
        RECT 396.955 -17.845 397.285 -17.515 ;
        RECT 395.595 -17.845 395.925 -17.515 ;
        RECT 392.875 -17.845 393.205 -17.515 ;
        RECT 391.515 -17.845 391.845 -17.515 ;
        RECT 390.155 -17.845 390.485 -17.515 ;
        RECT 388.795 -17.845 389.125 -17.515 ;
        RECT 387.435 -17.845 387.765 -17.515 ;
        RECT 386.075 -17.845 386.405 -17.515 ;
        RECT 384.715 -17.845 385.045 -17.515 ;
        RECT 383.355 -17.845 383.685 -17.515 ;
        RECT 381.995 -17.845 382.325 -17.515 ;
        RECT 380.635 -17.845 380.965 -17.515 ;
        RECT 377.915 -17.845 378.245 -17.515 ;
        RECT 376.555 -17.845 376.885 -17.515 ;
        RECT 375.195 -17.845 375.525 -17.515 ;
        RECT 373.835 -17.845 374.165 -17.515 ;
        RECT 372.475 -17.845 372.805 -17.515 ;
        RECT 371.115 -17.845 371.445 -17.515 ;
        RECT 369.755 -17.845 370.085 -17.515 ;
        RECT 368.395 -17.845 368.725 -17.515 ;
        RECT 367.035 -17.845 367.365 -17.515 ;
        RECT 365.675 -17.845 366.005 -17.515 ;
        RECT 362.955 -17.845 363.285 -17.515 ;
        RECT 361.595 -17.845 361.925 -17.515 ;
        RECT 360.235 -17.845 360.565 -17.515 ;
        RECT 358.875 -17.845 359.205 -17.515 ;
        RECT 357.515 -17.845 357.845 -17.515 ;
        RECT 356.155 -17.845 356.485 -17.515 ;
        RECT 354.795 -17.845 355.125 -17.515 ;
        RECT 353.435 -17.845 353.765 -17.515 ;
        RECT 352.075 -17.845 352.405 -17.515 ;
        RECT 350.715 -17.845 351.045 -17.515 ;
        RECT 347.995 -17.845 348.325 -17.515 ;
        RECT 346.635 -17.845 346.965 -17.515 ;
        RECT 345.275 -17.845 345.605 -17.515 ;
        RECT 343.915 -17.845 344.245 -17.515 ;
        RECT 342.555 -17.845 342.885 -17.515 ;
        RECT 341.195 -17.845 341.525 -17.515 ;
        RECT 339.835 -17.845 340.165 -17.515 ;
        RECT 338.475 -17.845 338.805 -17.515 ;
        RECT 337.115 -17.845 337.445 -17.515 ;
        RECT 335.755 -17.845 336.085 -17.515 ;
        RECT 333.035 -17.845 333.365 -17.515 ;
        RECT 331.675 -17.845 332.005 -17.515 ;
        RECT 330.315 -17.845 330.645 -17.515 ;
        RECT 328.955 -17.845 329.285 -17.515 ;
        RECT 327.595 -17.845 327.925 -17.515 ;
        RECT 326.235 -17.845 326.565 -17.515 ;
        RECT 324.875 -17.845 325.205 -17.515 ;
        RECT 323.515 -17.845 323.845 -17.515 ;
        RECT 322.155 -17.845 322.485 -17.515 ;
        RECT 320.795 -17.845 321.125 -17.515 ;
        RECT 318.075 -17.845 318.405 -17.515 ;
        RECT 316.715 -17.845 317.045 -17.515 ;
        RECT 315.355 -17.845 315.685 -17.515 ;
        RECT 313.995 -17.845 314.325 -17.515 ;
        RECT 312.635 -17.845 312.965 -17.515 ;
        RECT 311.275 -17.845 311.605 -17.515 ;
        RECT 309.915 -17.845 310.245 -17.515 ;
        RECT 308.555 -17.845 308.885 -17.515 ;
        RECT 307.195 -17.845 307.525 -17.515 ;
        RECT 305.835 -17.845 306.165 -17.515 ;
        RECT 303.115 -17.845 303.445 -17.515 ;
        RECT 301.755 -17.845 302.085 -17.515 ;
        RECT 300.395 -17.845 300.725 -17.515 ;
        RECT 299.035 -17.845 299.365 -17.515 ;
        RECT 297.675 -17.845 298.005 -17.515 ;
        RECT 296.315 -17.845 296.645 -17.515 ;
        RECT 294.955 -17.845 295.285 -17.515 ;
        RECT 293.595 -17.845 293.925 -17.515 ;
        RECT 292.235 -17.845 292.565 -17.515 ;
        RECT 290.875 -17.845 291.205 -17.515 ;
        RECT 288.155 -17.845 288.485 -17.515 ;
        RECT 286.795 -17.845 287.125 -17.515 ;
        RECT 285.435 -17.845 285.765 -17.515 ;
        RECT 284.075 -17.845 284.405 -17.515 ;
        RECT 282.715 -17.845 283.045 -17.515 ;
        RECT 281.355 -17.845 281.685 -17.515 ;
        RECT 279.995 -17.845 280.325 -17.515 ;
        RECT 278.635 -17.845 278.965 -17.515 ;
        RECT 277.275 -17.845 277.605 -17.515 ;
        RECT 275.915 -17.845 276.245 -17.515 ;
        RECT 273.195 -17.845 273.525 -17.515 ;
        RECT 271.835 -17.845 272.165 -17.515 ;
        RECT 270.475 -17.845 270.805 -17.515 ;
        RECT 269.115 -17.845 269.445 -17.515 ;
        RECT 267.755 -17.845 268.085 -17.515 ;
        RECT 266.395 -17.845 266.725 -17.515 ;
        RECT 265.035 -17.845 265.365 -17.515 ;
        RECT 263.675 -17.845 264.005 -17.515 ;
        RECT 262.315 -17.845 262.645 -17.515 ;
        RECT 260.955 -17.845 261.285 -17.515 ;
        RECT 258.235 -17.845 258.565 -17.515 ;
        RECT 256.875 -17.845 257.205 -17.515 ;
        RECT 255.515 -17.845 255.845 -17.515 ;
        RECT 254.155 -17.845 254.485 -17.515 ;
        RECT 252.795 -17.845 253.125 -17.515 ;
        RECT 251.435 -17.845 251.765 -17.515 ;
        RECT 250.075 -17.845 250.405 -17.515 ;
        RECT 248.715 -17.845 249.045 -17.515 ;
        RECT 247.355 -17.845 247.685 -17.515 ;
        RECT 245.995 -17.845 246.325 -17.515 ;
        RECT 243.275 -17.845 243.605 -17.515 ;
        RECT 241.915 -17.845 242.245 -17.515 ;
        RECT 240.555 -17.845 240.885 -17.515 ;
        RECT 239.195 -17.845 239.525 -17.515 ;
        RECT 237.835 -17.845 238.165 -17.515 ;
        RECT 236.475 -17.845 236.805 -17.515 ;
        RECT 235.115 -17.845 235.445 -17.515 ;
        RECT 233.755 -17.845 234.085 -17.515 ;
        RECT 232.395 -17.845 232.725 -17.515 ;
        RECT 231.035 -17.845 231.365 -17.515 ;
        RECT 228.315 -17.845 228.645 -17.515 ;
        RECT 226.955 -17.845 227.285 -17.515 ;
        RECT 225.595 -17.845 225.925 -17.515 ;
        RECT 224.235 -17.845 224.565 -17.515 ;
        RECT 222.875 -17.845 223.205 -17.515 ;
        RECT 221.515 -17.845 221.845 -17.515 ;
        RECT 220.155 -17.845 220.485 -17.515 ;
        RECT 218.795 -17.845 219.125 -17.515 ;
        RECT 217.435 -17.845 217.765 -17.515 ;
        RECT 216.075 -17.845 216.405 -17.515 ;
        RECT 213.355 -17.845 213.685 -17.515 ;
        RECT 211.995 -17.845 212.325 -17.515 ;
        RECT 210.635 -17.845 210.965 -17.515 ;
        RECT 209.275 -17.845 209.605 -17.515 ;
        RECT 207.915 -17.845 208.245 -17.515 ;
        RECT 206.555 -17.845 206.885 -17.515 ;
        RECT 205.195 -17.845 205.525 -17.515 ;
        RECT 203.835 -17.845 204.165 -17.515 ;
        RECT 202.475 -17.845 202.805 -17.515 ;
        RECT 201.115 -17.845 201.445 -17.515 ;
        RECT 198.395 -17.845 198.725 -17.515 ;
        RECT 197.035 -17.845 197.365 -17.515 ;
        RECT 195.675 -17.845 196.005 -17.515 ;
        RECT 194.315 -17.845 194.645 -17.515 ;
        RECT 192.955 -17.845 193.285 -17.515 ;
        RECT 191.595 -17.845 191.925 -17.515 ;
        RECT 190.235 -17.845 190.565 -17.515 ;
        RECT 188.875 -17.845 189.205 -17.515 ;
        RECT 187.515 -17.845 187.845 -17.515 ;
        RECT 186.155 -17.845 186.485 -17.515 ;
        RECT 183.435 -17.845 183.765 -17.515 ;
        RECT 182.075 -17.845 182.405 -17.515 ;
        RECT 180.715 -17.845 181.045 -17.515 ;
        RECT 179.355 -17.845 179.685 -17.515 ;
        RECT 177.995 -17.845 178.325 -17.515 ;
        RECT 176.635 -17.845 176.965 -17.515 ;
        RECT 175.275 -17.845 175.605 -17.515 ;
        RECT 173.915 -17.845 174.245 -17.515 ;
        RECT 172.555 -17.845 172.885 -17.515 ;
        RECT 171.195 -17.845 171.525 -17.515 ;
        RECT 168.475 -17.845 168.805 -17.515 ;
        RECT 167.115 -17.845 167.445 -17.515 ;
        RECT 165.755 -17.845 166.085 -17.515 ;
        RECT 164.395 -17.845 164.725 -17.515 ;
        RECT 163.035 -17.845 163.365 -17.515 ;
        RECT 161.675 -17.845 162.005 -17.515 ;
        RECT 160.315 -17.845 160.645 -17.515 ;
        RECT 158.955 -17.845 159.285 -17.515 ;
        RECT 157.595 -17.845 157.925 -17.515 ;
        RECT 156.235 -17.845 156.565 -17.515 ;
        RECT 153.515 -17.845 153.845 -17.515 ;
        RECT 152.155 -17.845 152.485 -17.515 ;
        RECT 150.795 -17.845 151.125 -17.515 ;
        RECT 149.435 -17.845 149.765 -17.515 ;
        RECT 148.075 -17.845 148.405 -17.515 ;
        RECT 146.715 -17.845 147.045 -17.515 ;
        RECT 145.355 -17.845 145.685 -17.515 ;
        RECT 143.995 -17.845 144.325 -17.515 ;
        RECT 142.635 -17.845 142.965 -17.515 ;
        RECT 141.275 -17.845 141.605 -17.515 ;
        RECT 138.555 -17.845 138.885 -17.515 ;
        RECT 137.195 -17.845 137.525 -17.515 ;
        RECT 135.835 -17.845 136.165 -17.515 ;
        RECT 134.475 -17.845 134.805 -17.515 ;
        RECT 133.115 -17.845 133.445 -17.515 ;
        RECT 131.755 -17.845 132.085 -17.515 ;
        RECT 130.395 -17.845 130.725 -17.515 ;
        RECT 129.035 -17.845 129.365 -17.515 ;
        RECT 127.675 -17.845 128.005 -17.515 ;
        RECT 126.315 -17.845 126.645 -17.515 ;
        RECT 123.595 -17.845 123.925 -17.515 ;
        RECT 122.235 -17.845 122.565 -17.515 ;
        RECT 120.875 -17.845 121.205 -17.515 ;
        RECT 119.515 -17.845 119.845 -17.515 ;
        RECT 118.155 -17.845 118.485 -17.515 ;
        RECT 116.795 -17.845 117.125 -17.515 ;
        RECT 115.435 -17.845 115.765 -17.515 ;
        RECT 114.075 -17.845 114.405 -17.515 ;
        RECT 112.715 -17.845 113.045 -17.515 ;
        RECT 111.355 -17.845 111.685 -17.515 ;
        RECT 108.635 -17.845 108.965 -17.515 ;
        RECT 107.275 -17.845 107.605 -17.515 ;
        RECT 105.915 -17.845 106.245 -17.515 ;
        RECT 104.555 -17.845 104.885 -17.515 ;
        RECT 103.195 -17.845 103.525 -17.515 ;
        RECT 101.835 -17.845 102.165 -17.515 ;
        RECT 100.475 -17.845 100.805 -17.515 ;
        RECT 99.115 -17.845 99.445 -17.515 ;
        RECT 97.755 -17.845 98.085 -17.515 ;
        RECT 96.395 -17.845 96.725 -17.515 ;
        RECT 93.675 -17.845 94.005 -17.515 ;
        RECT 92.315 -17.845 92.645 -17.515 ;
        RECT 90.955 -17.845 91.285 -17.515 ;
        RECT 89.595 -17.845 89.925 -17.515 ;
        RECT 88.235 -17.845 88.565 -17.515 ;
        RECT 86.875 -17.845 87.205 -17.515 ;
        RECT 85.515 -17.845 85.845 -17.515 ;
        RECT 84.155 -17.845 84.485 -17.515 ;
        RECT 82.795 -17.845 83.125 -17.515 ;
        RECT 81.435 -17.845 81.765 -17.515 ;
        RECT 80.075 -17.845 80.405 -17.515 ;
        RECT 78.715 -17.845 79.045 -17.515 ;
        RECT 77.355 -17.845 77.685 -17.515 ;
        RECT 75.995 -17.845 76.325 -17.515 ;
        RECT 74.635 -17.845 74.965 -17.515 ;
        RECT 73.275 -17.845 73.605 -17.515 ;
        RECT 71.915 -17.845 72.245 -17.515 ;
        RECT 70.555 -17.845 70.885 -17.515 ;
        RECT 69.195 -17.845 69.525 -17.515 ;
        RECT 67.835 -17.845 68.165 -17.515 ;
        RECT 65.115 -17.845 65.445 -17.515 ;
        RECT 63.755 -17.845 64.085 -17.515 ;
        RECT 62.395 -17.845 62.725 -17.515 ;
        RECT 61.035 -17.845 61.365 -17.515 ;
        RECT 59.675 -17.845 60.005 -17.515 ;
        RECT 58.315 -17.845 58.645 -17.515 ;
        RECT 56.955 -17.845 57.285 -17.515 ;
        RECT 55.595 -17.845 55.925 -17.515 ;
        RECT 54.235 -17.845 54.565 -17.515 ;
        RECT 52.875 -17.845 53.205 -17.515 ;
        RECT 50.155 -17.845 50.485 -17.515 ;
        RECT 48.795 -17.845 49.125 -17.515 ;
        RECT 47.435 -17.845 47.765 -17.515 ;
        RECT 46.075 -17.845 46.405 -17.515 ;
        RECT 44.715 -17.845 45.045 -17.515 ;
        RECT 43.355 -17.845 43.685 -17.515 ;
        RECT 41.995 -17.845 42.325 -17.515 ;
        RECT 40.635 -17.845 40.965 -17.515 ;
        RECT 39.275 -17.845 39.605 -17.515 ;
        RECT 37.915 -17.845 38.245 -17.515 ;
        RECT 35.195 -17.845 35.525 -17.515 ;
        RECT 33.835 -17.845 34.165 -17.515 ;
        RECT 32.475 -17.845 32.805 -17.515 ;
        RECT 31.115 -17.845 31.445 -17.515 ;
        RECT 29.755 -17.845 30.085 -17.515 ;
        RECT 28.395 -17.845 28.725 -17.515 ;
        RECT 27.035 -17.845 27.365 -17.515 ;
        RECT 25.675 -17.845 26.005 -17.515 ;
        RECT 24.315 -17.845 24.645 -17.515 ;
        RECT 22.955 -17.845 23.285 -17.515 ;
        RECT 20.235 -17.845 20.565 -17.515 ;
        RECT 18.875 -17.845 19.205 -17.515 ;
        RECT 17.515 -17.845 17.845 -17.515 ;
        RECT 16.155 -17.845 16.485 -17.515 ;
        RECT 14.795 -17.845 15.125 -17.515 ;
        RECT 13.435 -17.845 13.765 -17.515 ;
        RECT 12.075 -17.845 12.405 -17.515 ;
        RECT 10.715 -17.845 11.045 -17.515 ;
        RECT 9.355 -17.845 9.685 -17.515 ;
        RECT 7.995 -17.845 8.325 -17.515 ;
        RECT 6.635 -17.845 6.965 -17.515 ;
        RECT 5.275 -17.845 5.605 -17.515 ;
        RECT 3.915 -17.845 4.245 -17.515 ;
        RECT 2.555 -17.845 2.885 -17.515 ;
        RECT 1.195 -17.845 1.525 -17.515 ;
        RECT -0.165 -17.845 0.165 -17.515 ;
        RECT -1.525 -17.845 -1.195 -17.515 ;
        RECT 883.835 -17.845 884.165 -17.515 ;
        RECT 882.475 -17.845 882.805 -17.515 ;
        RECT 881.115 -17.845 881.445 -17.515 ;
        RECT 879.755 -17.845 880.085 -17.515 ;
        RECT 878.395 -17.845 878.725 -17.515 ;
        RECT 877.035 -17.845 877.365 -17.515 ;
        RECT 875.675 -17.845 876.005 -17.515 ;
        RECT 874.315 -17.845 874.645 -17.515 ;
        RECT 872.955 -17.845 873.285 -17.515 ;
        RECT 871.595 -17.845 871.925 -17.515 ;
        RECT 868.875 -17.845 869.205 -17.515 ;
        RECT 867.515 -17.845 867.845 -17.515 ;
        RECT 866.155 -17.845 866.485 -17.515 ;
        RECT 864.795 -17.845 865.125 -17.515 ;
        RECT 863.435 -17.845 863.765 -17.515 ;
        RECT 862.075 -17.845 862.405 -17.515 ;
        RECT 860.715 -17.845 861.045 -17.515 ;
        RECT 859.355 -17.845 859.685 -17.515 ;
        RECT 857.995 -17.845 858.325 -17.515 ;
        RECT 856.635 -17.845 856.965 -17.515 ;
        RECT 853.915 -17.845 854.245 -17.515 ;
        RECT 852.555 -17.845 852.885 -17.515 ;
        RECT 851.195 -17.845 851.525 -17.515 ;
        RECT 849.835 -17.845 850.165 -17.515 ;
        RECT 848.475 -17.845 848.805 -17.515 ;
        RECT 847.115 -17.845 847.445 -17.515 ;
        RECT 845.755 -17.845 846.085 -17.515 ;
        RECT 844.395 -17.845 844.725 -17.515 ;
        RECT 843.035 -17.845 843.365 -17.515 ;
        RECT 841.675 -17.845 842.005 -17.515 ;
        RECT 838.955 -17.845 839.285 -17.515 ;
        RECT 837.595 -17.845 837.925 -17.515 ;
        RECT 836.235 -17.845 836.565 -17.515 ;
        RECT 834.875 -17.845 835.205 -17.515 ;
        RECT 833.515 -17.845 833.845 -17.515 ;
        RECT 832.155 -17.845 832.485 -17.515 ;
        RECT 830.795 -17.845 831.125 -17.515 ;
        RECT 829.435 -17.845 829.765 -17.515 ;
        RECT 828.075 -17.845 828.405 -17.515 ;
        RECT 826.715 -17.845 827.045 -17.515 ;
        RECT 823.995 -17.845 824.325 -17.515 ;
        RECT 822.635 -17.845 822.965 -17.515 ;
        RECT 821.275 -17.845 821.605 -17.515 ;
        RECT 819.915 -17.845 820.245 -17.515 ;
        RECT 818.555 -17.845 818.885 -17.515 ;
        RECT 817.195 -17.845 817.525 -17.515 ;
        RECT 815.835 -17.845 816.165 -17.515 ;
        RECT 814.475 -17.845 814.805 -17.515 ;
        RECT 813.115 -17.845 813.445 -17.515 ;
        RECT 811.755 -17.845 812.085 -17.515 ;
        RECT 809.035 -17.845 809.365 -17.515 ;
        RECT 807.675 -17.845 808.005 -17.515 ;
        RECT 806.315 -17.845 806.645 -17.515 ;
        RECT 804.955 -17.845 805.285 -17.515 ;
        RECT 803.595 -17.845 803.925 -17.515 ;
        RECT 802.235 -17.845 802.565 -17.515 ;
        RECT 800.875 -17.845 801.205 -17.515 ;
        RECT 799.515 -17.845 799.845 -17.515 ;
        RECT 798.155 -17.845 798.485 -17.515 ;
        RECT 796.795 -17.845 797.125 -17.515 ;
        RECT 794.075 -17.845 794.405 -17.515 ;
        RECT 792.715 -17.845 793.045 -17.515 ;
        RECT 791.355 -17.845 791.685 -17.515 ;
        RECT 789.995 -17.845 790.325 -17.515 ;
        RECT 788.635 -17.845 788.965 -17.515 ;
        RECT 787.275 -17.845 787.605 -17.515 ;
        RECT 785.915 -17.845 786.245 -17.515 ;
        RECT 784.555 -17.845 784.885 -17.515 ;
        RECT 783.195 -17.845 783.525 -17.515 ;
        RECT 781.835 -17.845 782.165 -17.515 ;
        RECT 779.115 -17.845 779.445 -17.515 ;
        RECT 777.755 -17.845 778.085 -17.515 ;
        RECT 776.395 -17.845 776.725 -17.515 ;
        RECT 775.035 -17.845 775.365 -17.515 ;
        RECT 773.675 -17.845 774.005 -17.515 ;
        RECT 772.315 -17.845 772.645 -17.515 ;
        RECT 770.955 -17.845 771.285 -17.515 ;
        RECT 769.595 -17.845 769.925 -17.515 ;
        RECT 768.235 -17.845 768.565 -17.515 ;
        RECT 766.875 -17.845 767.205 -17.515 ;
        RECT 764.155 -17.845 764.485 -17.515 ;
        RECT 762.795 -17.845 763.125 -17.515 ;
        RECT 761.435 -17.845 761.765 -17.515 ;
        RECT 760.075 -17.845 760.405 -17.515 ;
        RECT 758.715 -17.845 759.045 -17.515 ;
        RECT 757.355 -17.845 757.685 -17.515 ;
        RECT 755.995 -17.845 756.325 -17.515 ;
        RECT 754.635 -17.845 754.965 -17.515 ;
        RECT 753.275 -17.845 753.605 -17.515 ;
        RECT 750.555 -17.845 750.885 -17.515 ;
        RECT 749.195 -17.845 749.525 -17.515 ;
        RECT 747.835 -17.845 748.165 -17.515 ;
        RECT 746.475 -17.845 746.805 -17.515 ;
        RECT 745.115 -17.845 745.445 -17.515 ;
        RECT 743.755 -17.845 744.085 -17.515 ;
        RECT 954.555 -17.845 954.885 -17.515 ;
        RECT 743.755 -17.84 954.885 -17.52 ;
        RECT 953.195 -17.845 953.525 -17.515 ;
        RECT 951.835 -17.845 952.165 -17.515 ;
        RECT 950.475 -17.845 950.805 -17.515 ;
        RECT 949.115 -17.845 949.445 -17.515 ;
        RECT 947.755 -17.845 948.085 -17.515 ;
        RECT 946.395 -17.845 946.725 -17.515 ;
        RECT 945.035 -17.845 945.365 -17.515 ;
        RECT 943.675 -17.845 944.005 -17.515 ;
        RECT 942.315 -17.845 942.645 -17.515 ;
        RECT 940.955 -17.845 941.285 -17.515 ;
        RECT 939.595 -17.845 939.925 -17.515 ;
        RECT 938.235 -17.845 938.565 -17.515 ;
        RECT 936.875 -17.845 937.205 -17.515 ;
        RECT 935.515 -17.845 935.845 -17.515 ;
        RECT 934.155 -17.845 934.485 -17.515 ;
        RECT 932.795 -17.845 933.125 -17.515 ;
        RECT 931.435 -17.845 931.765 -17.515 ;
        RECT 928.715 -17.845 929.045 -17.515 ;
        RECT 927.355 -17.845 927.685 -17.515 ;
        RECT 925.995 -17.845 926.325 -17.515 ;
        RECT 924.635 -17.845 924.965 -17.515 ;
        RECT 923.275 -17.845 923.605 -17.515 ;
        RECT 921.915 -17.845 922.245 -17.515 ;
        RECT 920.555 -17.845 920.885 -17.515 ;
        RECT 919.195 -17.845 919.525 -17.515 ;
        RECT 917.835 -17.845 918.165 -17.515 ;
        RECT 916.475 -17.845 916.805 -17.515 ;
        RECT 913.755 -17.845 914.085 -17.515 ;
        RECT 912.395 -17.845 912.725 -17.515 ;
        RECT 911.035 -17.845 911.365 -17.515 ;
        RECT 909.675 -17.845 910.005 -17.515 ;
        RECT 908.315 -17.845 908.645 -17.515 ;
        RECT 906.955 -17.845 907.285 -17.515 ;
        RECT 905.595 -17.845 905.925 -17.515 ;
        RECT 904.235 -17.845 904.565 -17.515 ;
        RECT 902.875 -17.845 903.205 -17.515 ;
        RECT 901.515 -17.845 901.845 -17.515 ;
        RECT 898.795 -17.845 899.125 -17.515 ;
        RECT 897.435 -17.845 897.765 -17.515 ;
        RECT 896.075 -17.845 896.405 -17.515 ;
        RECT 894.715 -17.845 895.045 -17.515 ;
        RECT 893.355 -17.845 893.685 -17.515 ;
        RECT 891.995 -17.845 892.325 -17.515 ;
        RECT 890.635 -17.845 890.965 -17.515 ;
        RECT 889.275 -17.845 889.605 -17.515 ;
        RECT 887.915 -17.845 888.245 -17.515 ;
        RECT 886.555 -17.845 886.885 -17.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.04 -30.08 747.48 -29.76 ;
        RECT 746.475 -30.085 746.805 -29.755 ;
        RECT 745.115 -30.085 745.445 -29.755 ;
        RECT 743.755 -30.085 744.085 -29.755 ;
        RECT 742.395 -30.085 742.725 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 736.96 -23.28 748.16 -22.96 ;
        RECT 746.475 -23.285 746.805 -22.955 ;
        RECT 745.115 -23.285 745.445 -22.955 ;
        RECT 743.755 -23.285 744.085 -22.955 ;
        RECT 742.395 -23.285 742.725 -22.955 ;
        RECT 741.035 -23.285 741.365 -22.955 ;
        RECT 738.315 -23.285 738.645 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 737.64 -27.36 748.16 -27.04 ;
        RECT 746.475 -27.365 746.805 -27.035 ;
        RECT 745.115 -27.365 745.445 -27.035 ;
        RECT 743.755 -27.365 744.085 -27.035 ;
        RECT 742.395 -27.365 742.725 -27.035 ;
        RECT 738.315 -27.365 738.645 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 747.835 -35.525 748.165 -35.195 ;
        RECT 741.04 -35.52 748.165 -35.2 ;
        RECT 746.475 -35.525 746.805 -35.195 ;
        RECT 745.115 -35.525 745.445 -35.195 ;
        RECT 743.755 -35.525 744.085 -35.195 ;
        RECT 742.395 -35.525 742.725 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 741.04 -26 751.56 -25.68 ;
        RECT 750.555 -26.005 750.885 -25.675 ;
        RECT 749.195 -26.005 749.525 -25.675 ;
        RECT 746.475 -26.005 746.805 -25.675 ;
        RECT 745.115 -26.005 745.445 -25.675 ;
        RECT 743.755 -26.005 744.085 -25.675 ;
        RECT 742.395 -26.005 742.725 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 756 -30.08 762.44 -29.76 ;
        RECT 761.435 -30.085 761.765 -29.755 ;
        RECT 760.075 -30.085 760.405 -29.755 ;
        RECT 758.715 -30.085 759.045 -29.755 ;
        RECT 757.355 -30.085 757.685 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 751.92 -23.28 763.12 -22.96 ;
        RECT 761.435 -23.285 761.765 -22.955 ;
        RECT 760.075 -23.285 760.405 -22.955 ;
        RECT 758.715 -23.285 759.045 -22.955 ;
        RECT 757.355 -23.285 757.685 -22.955 ;
        RECT 755.995 -23.285 756.325 -22.955 ;
        RECT 753.275 -23.285 753.605 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 752.6 -27.36 763.12 -27.04 ;
        RECT 761.435 -27.365 761.765 -27.035 ;
        RECT 760.075 -27.365 760.405 -27.035 ;
        RECT 758.715 -27.365 759.045 -27.035 ;
        RECT 757.355 -27.365 757.685 -27.035 ;
        RECT 753.275 -27.365 753.605 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 762.795 -35.525 763.125 -35.195 ;
        RECT 756 -35.52 763.125 -35.2 ;
        RECT 761.435 -35.525 761.765 -35.195 ;
        RECT 760.075 -35.525 760.405 -35.195 ;
        RECT 758.715 -35.525 759.045 -35.195 ;
        RECT 757.355 -35.525 757.685 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 756 -26 766.52 -25.68 ;
        RECT 764.155 -26.005 764.485 -25.675 ;
        RECT 761.435 -26.005 761.765 -25.675 ;
        RECT 760.075 -26.005 760.405 -25.675 ;
        RECT 758.715 -26.005 759.045 -25.675 ;
        RECT 757.355 -26.005 757.685 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 770.96 -30.08 777.4 -29.76 ;
        RECT 776.395 -30.085 776.725 -29.755 ;
        RECT 775.035 -30.085 775.365 -29.755 ;
        RECT 773.675 -30.085 774.005 -29.755 ;
        RECT 772.315 -30.085 772.645 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.875 -23.28 778.08 -22.96 ;
        RECT 776.395 -23.285 776.725 -22.955 ;
        RECT 775.035 -23.285 775.365 -22.955 ;
        RECT 773.675 -23.285 774.005 -22.955 ;
        RECT 772.315 -23.285 772.645 -22.955 ;
        RECT 770.955 -23.285 771.285 -22.955 ;
        RECT 768.235 -23.285 768.565 -22.955 ;
        RECT 766.875 -23.285 767.205 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 766.88 -27.36 778.08 -27.04 ;
        RECT 776.395 -27.365 776.725 -27.035 ;
        RECT 775.035 -27.365 775.365 -27.035 ;
        RECT 773.675 -27.365 774.005 -27.035 ;
        RECT 772.315 -27.365 772.645 -27.035 ;
        RECT 768.235 -27.365 768.565 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 777.755 -35.525 778.085 -35.195 ;
        RECT 770.96 -35.52 778.085 -35.2 ;
        RECT 776.395 -35.525 776.725 -35.195 ;
        RECT 775.035 -35.525 775.365 -35.195 ;
        RECT 773.675 -35.525 774.005 -35.195 ;
        RECT 772.315 -35.525 772.645 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 770.96 -26 781.48 -25.68 ;
        RECT 779.115 -26.005 779.445 -25.675 ;
        RECT 776.395 -26.005 776.725 -25.675 ;
        RECT 775.035 -26.005 775.365 -25.675 ;
        RECT 773.675 -26.005 774.005 -25.675 ;
        RECT 772.315 -26.005 772.645 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 785.92 -30.08 792.36 -29.76 ;
        RECT 791.355 -30.085 791.685 -29.755 ;
        RECT 789.995 -30.085 790.325 -29.755 ;
        RECT 788.635 -30.085 788.965 -29.755 ;
        RECT 787.275 -30.085 787.605 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 781.16 -23.28 793.04 -22.96 ;
        RECT 791.355 -23.285 791.685 -22.955 ;
        RECT 789.995 -23.285 790.325 -22.955 ;
        RECT 788.635 -23.285 788.965 -22.955 ;
        RECT 787.275 -23.285 787.605 -22.955 ;
        RECT 785.915 -23.285 786.245 -22.955 ;
        RECT 783.195 -23.285 783.525 -22.955 ;
        RECT 781.835 -23.285 782.165 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 781.84 -27.36 793.04 -27.04 ;
        RECT 791.355 -27.365 791.685 -27.035 ;
        RECT 789.995 -27.365 790.325 -27.035 ;
        RECT 788.635 -27.365 788.965 -27.035 ;
        RECT 787.275 -27.365 787.605 -27.035 ;
        RECT 783.195 -27.365 783.525 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 792.715 -35.525 793.045 -35.195 ;
        RECT 785.92 -35.52 793.045 -35.2 ;
        RECT 791.355 -35.525 791.685 -35.195 ;
        RECT 789.995 -35.525 790.325 -35.195 ;
        RECT 788.635 -35.525 788.965 -35.195 ;
        RECT 787.275 -35.525 787.605 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 785.92 -26 796.44 -25.68 ;
        RECT 794.075 -26.005 794.405 -25.675 ;
        RECT 791.355 -26.005 791.685 -25.675 ;
        RECT 789.995 -26.005 790.325 -25.675 ;
        RECT 788.635 -26.005 788.965 -25.675 ;
        RECT 787.275 -26.005 787.605 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 796.12 -23.28 807.32 -22.96 ;
        RECT 804.955 -23.285 805.285 -22.955 ;
        RECT 803.595 -23.285 803.925 -22.955 ;
        RECT 802.235 -23.285 802.565 -22.955 ;
        RECT 800.875 -23.285 801.205 -22.955 ;
        RECT 798.155 -23.285 798.485 -22.955 ;
        RECT 796.795 -23.285 797.125 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 796.8 -27.36 807.32 -27.04 ;
        RECT 804.955 -27.365 805.285 -27.035 ;
        RECT 803.595 -27.365 803.925 -27.035 ;
        RECT 802.235 -27.365 802.565 -27.035 ;
        RECT 798.155 -27.365 798.485 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 800.88 -30.08 807.32 -29.76 ;
        RECT 804.955 -30.085 805.285 -29.755 ;
        RECT 803.595 -30.085 803.925 -29.755 ;
        RECT 802.235 -30.085 802.565 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 800.88 -35.52 807.32 -35.2 ;
        RECT 806.315 -35.525 806.645 -35.195 ;
        RECT 804.955 -35.525 805.285 -35.195 ;
        RECT 803.595 -35.525 803.925 -35.195 ;
        RECT 802.235 -35.525 802.565 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 800.88 -26 811.4 -25.68 ;
        RECT 809.035 -26.005 809.365 -25.675 ;
        RECT 804.955 -26.005 805.285 -25.675 ;
        RECT 803.595 -26.005 803.925 -25.675 ;
        RECT 802.235 -26.005 802.565 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 815.84 -30.08 821.6 -29.76 ;
        RECT 819.915 -30.085 820.245 -29.755 ;
        RECT 818.555 -30.085 818.885 -29.755 ;
        RECT 817.195 -30.085 817.525 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 811.08 -23.28 822.28 -22.96 ;
        RECT 819.915 -23.285 820.245 -22.955 ;
        RECT 818.555 -23.285 818.885 -22.955 ;
        RECT 817.195 -23.285 817.525 -22.955 ;
        RECT 815.835 -23.285 816.165 -22.955 ;
        RECT 813.115 -23.285 813.445 -22.955 ;
        RECT 811.755 -23.285 812.085 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 811.76 -27.36 822.28 -27.04 ;
        RECT 819.915 -27.365 820.245 -27.035 ;
        RECT 818.555 -27.365 818.885 -27.035 ;
        RECT 817.195 -27.365 817.525 -27.035 ;
        RECT 813.115 -27.365 813.445 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 815.84 -35.52 822.28 -35.2 ;
        RECT 821.275 -35.525 821.605 -35.195 ;
        RECT 819.915 -35.525 820.245 -35.195 ;
        RECT 818.555 -35.525 818.885 -35.195 ;
        RECT 817.195 -35.525 817.525 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 815.84 -26 826.36 -25.68 ;
        RECT 823.995 -26.005 824.325 -25.675 ;
        RECT 819.915 -26.005 820.245 -25.675 ;
        RECT 818.555 -26.005 818.885 -25.675 ;
        RECT 817.195 -26.005 817.525 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 830.8 -30.08 836.56 -29.76 ;
        RECT 834.875 -30.085 835.205 -29.755 ;
        RECT 833.515 -30.085 833.845 -29.755 ;
        RECT 832.155 -30.085 832.485 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 826.04 -23.28 837.24 -22.96 ;
        RECT 834.875 -23.285 835.205 -22.955 ;
        RECT 833.515 -23.285 833.845 -22.955 ;
        RECT 832.155 -23.285 832.485 -22.955 ;
        RECT 830.795 -23.285 831.125 -22.955 ;
        RECT 828.075 -23.285 828.405 -22.955 ;
        RECT 826.715 -23.285 827.045 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 826.72 -27.36 837.24 -27.04 ;
        RECT 834.875 -27.365 835.205 -27.035 ;
        RECT 833.515 -27.365 833.845 -27.035 ;
        RECT 832.155 -27.365 832.485 -27.035 ;
        RECT 828.075 -27.365 828.405 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 830.8 -35.52 837.24 -35.2 ;
        RECT 836.235 -35.525 836.565 -35.195 ;
        RECT 834.875 -35.525 835.205 -35.195 ;
        RECT 833.515 -35.525 833.845 -35.195 ;
        RECT 832.155 -35.525 832.485 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 830.8 -26 841.32 -25.68 ;
        RECT 838.955 -26.005 839.285 -25.675 ;
        RECT 834.875 -26.005 835.205 -25.675 ;
        RECT 833.515 -26.005 833.845 -25.675 ;
        RECT 832.155 -26.005 832.485 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 845.755 -30.08 851.52 -29.76 ;
        RECT 849.835 -30.085 850.165 -29.755 ;
        RECT 848.475 -30.085 848.805 -29.755 ;
        RECT 847.115 -30.085 847.445 -29.755 ;
        RECT 845.755 -30.085 846.085 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 841 -23.28 852.2 -22.96 ;
        RECT 849.835 -23.285 850.165 -22.955 ;
        RECT 848.475 -23.285 848.805 -22.955 ;
        RECT 847.115 -23.285 847.445 -22.955 ;
        RECT 845.755 -23.285 846.085 -22.955 ;
        RECT 843.035 -23.285 843.365 -22.955 ;
        RECT 841.675 -23.285 842.005 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 841.68 -27.36 852.2 -27.04 ;
        RECT 849.835 -27.365 850.165 -27.035 ;
        RECT 848.475 -27.365 848.805 -27.035 ;
        RECT 847.115 -27.365 847.445 -27.035 ;
        RECT 845.755 -27.365 846.085 -27.035 ;
        RECT 843.035 -27.365 843.365 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 845.755 -35.52 852.2 -35.2 ;
        RECT 851.195 -35.525 851.525 -35.195 ;
        RECT 849.835 -35.525 850.165 -35.195 ;
        RECT 848.475 -35.525 848.805 -35.195 ;
        RECT 847.115 -35.525 847.445 -35.195 ;
        RECT 845.755 -35.525 846.085 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 845.755 -26 856.28 -25.68 ;
        RECT 853.915 -26.005 854.245 -25.675 ;
        RECT 849.835 -26.005 850.165 -25.675 ;
        RECT 848.475 -26.005 848.805 -25.675 ;
        RECT 847.115 -26.005 847.445 -25.675 ;
        RECT 845.755 -26.005 846.085 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 860.04 -30.08 866.48 -29.76 ;
        RECT 864.795 -30.085 865.125 -29.755 ;
        RECT 863.435 -30.085 863.765 -29.755 ;
        RECT 862.075 -30.085 862.405 -29.755 ;
        RECT 860.715 -30.085 861.045 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 855.96 -23.28 867.16 -22.96 ;
        RECT 864.795 -23.285 865.125 -22.955 ;
        RECT 863.435 -23.285 863.765 -22.955 ;
        RECT 862.075 -23.285 862.405 -22.955 ;
        RECT 860.715 -23.285 861.045 -22.955 ;
        RECT 857.995 -23.285 858.325 -22.955 ;
        RECT 856.635 -23.285 856.965 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 856.64 -27.36 867.16 -27.04 ;
        RECT 864.795 -27.365 865.125 -27.035 ;
        RECT 863.435 -27.365 863.765 -27.035 ;
        RECT 862.075 -27.365 862.405 -27.035 ;
        RECT 860.715 -27.365 861.045 -27.035 ;
        RECT 857.995 -27.365 858.325 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 860.04 -35.52 867.16 -35.2 ;
        RECT 866.155 -35.525 866.485 -35.195 ;
        RECT 864.795 -35.525 865.125 -35.195 ;
        RECT 863.435 -35.525 863.765 -35.195 ;
        RECT 862.075 -35.525 862.405 -35.195 ;
        RECT 860.715 -35.525 861.045 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 860.04 -26 871.24 -25.68 ;
        RECT 868.875 -26.005 869.205 -25.675 ;
        RECT 864.795 -26.005 865.125 -25.675 ;
        RECT 863.435 -26.005 863.765 -25.675 ;
        RECT 862.075 -26.005 862.405 -25.675 ;
        RECT 860.715 -26.005 861.045 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 875 -30.08 881.44 -29.76 ;
        RECT 879.755 -30.085 880.085 -29.755 ;
        RECT 878.395 -30.085 878.725 -29.755 ;
        RECT 877.035 -30.085 877.365 -29.755 ;
        RECT 875.675 -30.085 876.005 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 870.92 -23.28 882.12 -22.96 ;
        RECT 879.755 -23.285 880.085 -22.955 ;
        RECT 878.395 -23.285 878.725 -22.955 ;
        RECT 877.035 -23.285 877.365 -22.955 ;
        RECT 875.675 -23.285 876.005 -22.955 ;
        RECT 871.595 -23.285 871.925 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 871.6 -27.36 882.12 -27.04 ;
        RECT 879.755 -27.365 880.085 -27.035 ;
        RECT 878.395 -27.365 878.725 -27.035 ;
        RECT 877.035 -27.365 877.365 -27.035 ;
        RECT 875.675 -27.365 876.005 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 875 -35.52 882.12 -35.2 ;
        RECT 881.115 -35.525 881.445 -35.195 ;
        RECT 879.755 -35.525 880.085 -35.195 ;
        RECT 878.395 -35.525 878.725 -35.195 ;
        RECT 877.035 -35.525 877.365 -35.195 ;
        RECT 875.675 -35.525 876.005 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 875 -26 886.2 -25.68 ;
        RECT 883.835 -26.005 884.165 -25.675 ;
        RECT 879.755 -26.005 880.085 -25.675 ;
        RECT 878.395 -26.005 878.725 -25.675 ;
        RECT 877.035 -26.005 877.365 -25.675 ;
        RECT 875.675 -26.005 876.005 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 889.96 -30.08 896.4 -29.76 ;
        RECT 894.715 -30.085 895.045 -29.755 ;
        RECT 893.355 -30.085 893.685 -29.755 ;
        RECT 891.995 -30.085 892.325 -29.755 ;
        RECT 890.635 -30.085 890.965 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 885.88 -23.28 897.08 -22.96 ;
        RECT 894.715 -23.285 895.045 -22.955 ;
        RECT 893.355 -23.285 893.685 -22.955 ;
        RECT 891.995 -23.285 892.325 -22.955 ;
        RECT 890.635 -23.285 890.965 -22.955 ;
        RECT 886.555 -23.285 886.885 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 886.56 -27.36 897.08 -27.04 ;
        RECT 894.715 -27.365 895.045 -27.035 ;
        RECT 893.355 -27.365 893.685 -27.035 ;
        RECT 891.995 -27.365 892.325 -27.035 ;
        RECT 890.635 -27.365 890.965 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 889.96 -35.52 897.08 -35.2 ;
        RECT 896.075 -35.525 896.405 -35.195 ;
        RECT 894.715 -35.525 895.045 -35.195 ;
        RECT 893.355 -35.525 893.685 -35.195 ;
        RECT 891.995 -35.525 892.325 -35.195 ;
        RECT 890.635 -35.525 890.965 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 889.96 -26 900.48 -25.68 ;
        RECT 898.795 -26.005 899.125 -25.675 ;
        RECT 894.715 -26.005 895.045 -25.675 ;
        RECT 893.355 -26.005 893.685 -25.675 ;
        RECT 891.995 -26.005 892.325 -25.675 ;
        RECT 890.635 -26.005 890.965 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 904.92 -30.08 911.36 -29.76 ;
        RECT 909.675 -30.085 910.005 -29.755 ;
        RECT 908.315 -30.085 908.645 -29.755 ;
        RECT 906.955 -30.085 907.285 -29.755 ;
        RECT 905.595 -30.085 905.925 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 900.84 -23.28 912.04 -22.96 ;
        RECT 909.675 -23.285 910.005 -22.955 ;
        RECT 908.315 -23.285 908.645 -22.955 ;
        RECT 906.955 -23.285 907.285 -22.955 ;
        RECT 905.595 -23.285 905.925 -22.955 ;
        RECT 901.515 -23.285 901.845 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 901.52 -27.36 912.04 -27.04 ;
        RECT 909.675 -27.365 910.005 -27.035 ;
        RECT 908.315 -27.365 908.645 -27.035 ;
        RECT 906.955 -27.365 907.285 -27.035 ;
        RECT 905.595 -27.365 905.925 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 904.92 -35.52 912.04 -35.2 ;
        RECT 911.035 -35.525 911.365 -35.195 ;
        RECT 909.675 -35.525 910.005 -35.195 ;
        RECT 908.315 -35.525 908.645 -35.195 ;
        RECT 906.955 -35.525 907.285 -35.195 ;
        RECT 905.595 -35.525 905.925 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 904.92 -26 915.44 -25.68 ;
        RECT 913.755 -26.005 914.085 -25.675 ;
        RECT 909.675 -26.005 910.005 -25.675 ;
        RECT 908.315 -26.005 908.645 -25.675 ;
        RECT 906.955 -26.005 907.285 -25.675 ;
        RECT 905.595 -26.005 905.925 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -19.205 11.045 -18.875 ;
        RECT 9.355 -19.205 9.685 -18.875 ;
        RECT 7.995 -19.205 8.325 -18.875 ;
        RECT 6.635 -19.205 6.965 -18.875 ;
        RECT 3.915 -19.205 4.245 -18.875 ;
        RECT 2.555 -19.205 2.885 -18.875 ;
        RECT 1.195 -19.205 1.525 -18.875 ;
        RECT -0.165 -19.205 0.165 -18.875 ;
        RECT -1.525 -19.205 -1.195 -18.875 ;
        RECT -1.525 -19.2 920.555 -18.88 ;
        RECT 919.195 -19.205 919.525 -18.875 ;
        RECT 917.835 -19.205 918.165 -18.875 ;
        RECT 916.475 -19.205 916.805 -18.875 ;
        RECT 911.035 -19.205 911.365 -18.875 ;
        RECT 909.675 -19.205 910.005 -18.875 ;
        RECT 908.315 -19.205 908.645 -18.875 ;
        RECT 906.955 -19.205 907.285 -18.875 ;
        RECT 905.595 -19.205 905.925 -18.875 ;
        RECT 904.235 -19.205 904.565 -18.875 ;
        RECT 902.875 -19.205 903.205 -18.875 ;
        RECT 901.515 -19.205 901.845 -18.875 ;
        RECT 896.075 -19.205 896.405 -18.875 ;
        RECT 894.715 -19.205 895.045 -18.875 ;
        RECT 893.355 -19.205 893.685 -18.875 ;
        RECT 891.995 -19.205 892.325 -18.875 ;
        RECT 890.635 -19.205 890.965 -18.875 ;
        RECT 889.275 -19.205 889.605 -18.875 ;
        RECT 887.915 -19.205 888.245 -18.875 ;
        RECT 886.555 -19.205 886.885 -18.875 ;
        RECT 881.115 -19.205 881.445 -18.875 ;
        RECT 879.755 -19.205 880.085 -18.875 ;
        RECT 878.395 -19.205 878.725 -18.875 ;
        RECT 877.035 -19.205 877.365 -18.875 ;
        RECT 875.675 -19.205 876.005 -18.875 ;
        RECT 874.315 -19.205 874.645 -18.875 ;
        RECT 872.955 -19.205 873.285 -18.875 ;
        RECT 871.595 -19.205 871.925 -18.875 ;
        RECT 866.155 -19.205 866.485 -18.875 ;
        RECT 864.795 -19.205 865.125 -18.875 ;
        RECT 863.435 -19.205 863.765 -18.875 ;
        RECT 862.075 -19.205 862.405 -18.875 ;
        RECT 860.715 -19.205 861.045 -18.875 ;
        RECT 859.355 -19.205 859.685 -18.875 ;
        RECT 857.995 -19.205 858.325 -18.875 ;
        RECT 856.635 -19.205 856.965 -18.875 ;
        RECT 851.195 -19.205 851.525 -18.875 ;
        RECT 849.835 -19.205 850.165 -18.875 ;
        RECT 848.475 -19.205 848.805 -18.875 ;
        RECT 847.115 -19.205 847.445 -18.875 ;
        RECT 845.755 -19.205 846.085 -18.875 ;
        RECT 844.395 -19.205 844.725 -18.875 ;
        RECT 843.035 -19.205 843.365 -18.875 ;
        RECT 841.675 -19.205 842.005 -18.875 ;
        RECT 836.235 -19.205 836.565 -18.875 ;
        RECT 834.875 -19.205 835.205 -18.875 ;
        RECT 833.515 -19.205 833.845 -18.875 ;
        RECT 832.155 -19.205 832.485 -18.875 ;
        RECT 830.795 -19.205 831.125 -18.875 ;
        RECT 829.435 -19.205 829.765 -18.875 ;
        RECT 828.075 -19.205 828.405 -18.875 ;
        RECT 826.715 -19.205 827.045 -18.875 ;
        RECT 821.275 -19.205 821.605 -18.875 ;
        RECT 819.915 -19.205 820.245 -18.875 ;
        RECT 818.555 -19.205 818.885 -18.875 ;
        RECT 817.195 -19.205 817.525 -18.875 ;
        RECT 815.835 -19.205 816.165 -18.875 ;
        RECT 814.475 -19.205 814.805 -18.875 ;
        RECT 813.115 -19.205 813.445 -18.875 ;
        RECT 811.755 -19.205 812.085 -18.875 ;
        RECT 806.315 -19.205 806.645 -18.875 ;
        RECT 804.955 -19.205 805.285 -18.875 ;
        RECT 803.595 -19.205 803.925 -18.875 ;
        RECT 802.235 -19.205 802.565 -18.875 ;
        RECT 800.875 -19.205 801.205 -18.875 ;
        RECT 799.515 -19.205 799.845 -18.875 ;
        RECT 798.155 -19.205 798.485 -18.875 ;
        RECT 796.795 -19.205 797.125 -18.875 ;
        RECT 791.355 -19.205 791.685 -18.875 ;
        RECT 789.995 -19.205 790.325 -18.875 ;
        RECT 788.635 -19.205 788.965 -18.875 ;
        RECT 787.275 -19.205 787.605 -18.875 ;
        RECT 785.915 -19.205 786.245 -18.875 ;
        RECT 784.555 -19.205 784.885 -18.875 ;
        RECT 783.195 -19.205 783.525 -18.875 ;
        RECT 781.835 -19.205 782.165 -18.875 ;
        RECT 779.115 -19.205 779.445 -18.875 ;
        RECT 776.395 -19.205 776.725 -18.875 ;
        RECT 775.035 -19.205 775.365 -18.875 ;
        RECT 773.675 -19.205 774.005 -18.875 ;
        RECT 772.315 -19.205 772.645 -18.875 ;
        RECT 770.955 -19.205 771.285 -18.875 ;
        RECT 769.595 -19.205 769.925 -18.875 ;
        RECT 768.235 -19.205 768.565 -18.875 ;
        RECT 766.875 -19.205 767.205 -18.875 ;
        RECT 764.155 -19.205 764.485 -18.875 ;
        RECT 761.435 -19.205 761.765 -18.875 ;
        RECT 760.075 -19.205 760.405 -18.875 ;
        RECT 758.715 -19.205 759.045 -18.875 ;
        RECT 757.355 -19.205 757.685 -18.875 ;
        RECT 755.995 -19.205 756.325 -18.875 ;
        RECT 754.635 -19.205 754.965 -18.875 ;
        RECT 753.275 -19.205 753.605 -18.875 ;
        RECT 749.195 -19.205 749.525 -18.875 ;
        RECT 746.475 -19.205 746.805 -18.875 ;
        RECT 745.115 -19.205 745.445 -18.875 ;
        RECT 743.755 -19.205 744.085 -18.875 ;
        RECT 742.395 -19.205 742.725 -18.875 ;
        RECT 741.035 -19.205 741.365 -18.875 ;
        RECT 739.675 -19.205 740.005 -18.875 ;
        RECT 738.315 -19.205 738.645 -18.875 ;
        RECT 734.235 -19.205 734.565 -18.875 ;
        RECT 731.515 -19.205 731.845 -18.875 ;
        RECT 730.155 -19.205 730.485 -18.875 ;
        RECT 728.795 -19.205 729.125 -18.875 ;
        RECT 727.435 -19.205 727.765 -18.875 ;
        RECT 726.075 -19.205 726.405 -18.875 ;
        RECT 724.715 -19.205 725.045 -18.875 ;
        RECT 723.355 -19.205 723.685 -18.875 ;
        RECT 719.275 -19.205 719.605 -18.875 ;
        RECT 716.555 -19.205 716.885 -18.875 ;
        RECT 715.195 -19.205 715.525 -18.875 ;
        RECT 713.835 -19.205 714.165 -18.875 ;
        RECT 712.475 -19.205 712.805 -18.875 ;
        RECT 711.115 -19.205 711.445 -18.875 ;
        RECT 709.755 -19.205 710.085 -18.875 ;
        RECT 708.395 -19.205 708.725 -18.875 ;
        RECT 704.315 -19.205 704.645 -18.875 ;
        RECT 701.595 -19.205 701.925 -18.875 ;
        RECT 700.235 -19.205 700.565 -18.875 ;
        RECT 698.875 -19.205 699.205 -18.875 ;
        RECT 697.515 -19.205 697.845 -18.875 ;
        RECT 696.155 -19.205 696.485 -18.875 ;
        RECT 694.795 -19.205 695.125 -18.875 ;
        RECT 693.435 -19.205 693.765 -18.875 ;
        RECT 689.355 -19.205 689.685 -18.875 ;
        RECT 686.635 -19.205 686.965 -18.875 ;
        RECT 685.275 -19.205 685.605 -18.875 ;
        RECT 683.915 -19.205 684.245 -18.875 ;
        RECT 682.555 -19.205 682.885 -18.875 ;
        RECT 681.195 -19.205 681.525 -18.875 ;
        RECT 679.835 -19.205 680.165 -18.875 ;
        RECT 678.475 -19.205 678.805 -18.875 ;
        RECT 674.395 -19.205 674.725 -18.875 ;
        RECT 671.675 -19.205 672.005 -18.875 ;
        RECT 670.315 -19.205 670.645 -18.875 ;
        RECT 668.955 -19.205 669.285 -18.875 ;
        RECT 667.595 -19.205 667.925 -18.875 ;
        RECT 666.235 -19.205 666.565 -18.875 ;
        RECT 664.875 -19.205 665.205 -18.875 ;
        RECT 663.515 -19.205 663.845 -18.875 ;
        RECT 659.435 -19.205 659.765 -18.875 ;
        RECT 656.715 -19.205 657.045 -18.875 ;
        RECT 655.355 -19.205 655.685 -18.875 ;
        RECT 653.995 -19.205 654.325 -18.875 ;
        RECT 652.635 -19.205 652.965 -18.875 ;
        RECT 651.275 -19.205 651.605 -18.875 ;
        RECT 649.915 -19.205 650.245 -18.875 ;
        RECT 648.555 -19.205 648.885 -18.875 ;
        RECT 643.115 -19.205 643.445 -18.875 ;
        RECT 641.755 -19.205 642.085 -18.875 ;
        RECT 640.395 -19.205 640.725 -18.875 ;
        RECT 639.035 -19.205 639.365 -18.875 ;
        RECT 637.675 -19.205 638.005 -18.875 ;
        RECT 636.315 -19.205 636.645 -18.875 ;
        RECT 634.955 -19.205 635.285 -18.875 ;
        RECT 633.595 -19.205 633.925 -18.875 ;
        RECT 628.155 -19.205 628.485 -18.875 ;
        RECT 626.795 -19.205 627.125 -18.875 ;
        RECT 625.435 -19.205 625.765 -18.875 ;
        RECT 624.075 -19.205 624.405 -18.875 ;
        RECT 622.715 -19.205 623.045 -18.875 ;
        RECT 621.355 -19.205 621.685 -18.875 ;
        RECT 619.995 -19.205 620.325 -18.875 ;
        RECT 618.635 -19.205 618.965 -18.875 ;
        RECT 613.195 -19.205 613.525 -18.875 ;
        RECT 611.835 -19.205 612.165 -18.875 ;
        RECT 610.475 -19.205 610.805 -18.875 ;
        RECT 609.115 -19.205 609.445 -18.875 ;
        RECT 607.755 -19.205 608.085 -18.875 ;
        RECT 606.395 -19.205 606.725 -18.875 ;
        RECT 605.035 -19.205 605.365 -18.875 ;
        RECT 603.675 -19.205 604.005 -18.875 ;
        RECT 598.235 -19.205 598.565 -18.875 ;
        RECT 596.875 -19.205 597.205 -18.875 ;
        RECT 595.515 -19.205 595.845 -18.875 ;
        RECT 594.155 -19.205 594.485 -18.875 ;
        RECT 592.795 -19.205 593.125 -18.875 ;
        RECT 591.435 -19.205 591.765 -18.875 ;
        RECT 590.075 -19.205 590.405 -18.875 ;
        RECT 588.715 -19.205 589.045 -18.875 ;
        RECT 583.275 -19.205 583.605 -18.875 ;
        RECT 581.915 -19.205 582.245 -18.875 ;
        RECT 580.555 -19.205 580.885 -18.875 ;
        RECT 579.195 -19.205 579.525 -18.875 ;
        RECT 577.835 -19.205 578.165 -18.875 ;
        RECT 576.475 -19.205 576.805 -18.875 ;
        RECT 575.115 -19.205 575.445 -18.875 ;
        RECT 573.755 -19.205 574.085 -18.875 ;
        RECT 568.315 -19.205 568.645 -18.875 ;
        RECT 566.955 -19.205 567.285 -18.875 ;
        RECT 565.595 -19.205 565.925 -18.875 ;
        RECT 564.235 -19.205 564.565 -18.875 ;
        RECT 562.875 -19.205 563.205 -18.875 ;
        RECT 561.515 -19.205 561.845 -18.875 ;
        RECT 560.155 -19.205 560.485 -18.875 ;
        RECT 558.795 -19.205 559.125 -18.875 ;
        RECT 553.355 -19.205 553.685 -18.875 ;
        RECT 551.995 -19.205 552.325 -18.875 ;
        RECT 550.635 -19.205 550.965 -18.875 ;
        RECT 549.275 -19.205 549.605 -18.875 ;
        RECT 547.915 -19.205 548.245 -18.875 ;
        RECT 546.555 -19.205 546.885 -18.875 ;
        RECT 545.195 -19.205 545.525 -18.875 ;
        RECT 543.835 -19.205 544.165 -18.875 ;
        RECT 538.395 -19.205 538.725 -18.875 ;
        RECT 537.035 -19.205 537.365 -18.875 ;
        RECT 535.675 -19.205 536.005 -18.875 ;
        RECT 534.315 -19.205 534.645 -18.875 ;
        RECT 532.955 -19.205 533.285 -18.875 ;
        RECT 531.595 -19.205 531.925 -18.875 ;
        RECT 530.235 -19.205 530.565 -18.875 ;
        RECT 528.875 -19.205 529.205 -18.875 ;
        RECT 523.435 -19.205 523.765 -18.875 ;
        RECT 522.075 -19.205 522.405 -18.875 ;
        RECT 520.715 -19.205 521.045 -18.875 ;
        RECT 519.355 -19.205 519.685 -18.875 ;
        RECT 517.995 -19.205 518.325 -18.875 ;
        RECT 516.635 -19.205 516.965 -18.875 ;
        RECT 515.275 -19.205 515.605 -18.875 ;
        RECT 513.915 -19.205 514.245 -18.875 ;
        RECT 508.475 -19.205 508.805 -18.875 ;
        RECT 507.115 -19.205 507.445 -18.875 ;
        RECT 505.755 -19.205 506.085 -18.875 ;
        RECT 504.395 -19.205 504.725 -18.875 ;
        RECT 503.035 -19.205 503.365 -18.875 ;
        RECT 501.675 -19.205 502.005 -18.875 ;
        RECT 500.315 -19.205 500.645 -18.875 ;
        RECT 498.955 -19.205 499.285 -18.875 ;
        RECT 493.515 -19.205 493.845 -18.875 ;
        RECT 492.155 -19.205 492.485 -18.875 ;
        RECT 490.795 -19.205 491.125 -18.875 ;
        RECT 489.435 -19.205 489.765 -18.875 ;
        RECT 488.075 -19.205 488.405 -18.875 ;
        RECT 486.715 -19.205 487.045 -18.875 ;
        RECT 485.355 -19.205 485.685 -18.875 ;
        RECT 483.995 -19.205 484.325 -18.875 ;
        RECT 478.555 -19.205 478.885 -18.875 ;
        RECT 477.195 -19.205 477.525 -18.875 ;
        RECT 475.835 -19.205 476.165 -18.875 ;
        RECT 474.475 -19.205 474.805 -18.875 ;
        RECT 473.115 -19.205 473.445 -18.875 ;
        RECT 471.755 -19.205 472.085 -18.875 ;
        RECT 470.395 -19.205 470.725 -18.875 ;
        RECT 469.035 -19.205 469.365 -18.875 ;
        RECT 463.595 -19.205 463.925 -18.875 ;
        RECT 462.235 -19.205 462.565 -18.875 ;
        RECT 460.875 -19.205 461.205 -18.875 ;
        RECT 459.515 -19.205 459.845 -18.875 ;
        RECT 458.155 -19.205 458.485 -18.875 ;
        RECT 456.795 -19.205 457.125 -18.875 ;
        RECT 455.435 -19.205 455.765 -18.875 ;
        RECT 454.075 -19.205 454.405 -18.875 ;
        RECT 448.635 -19.205 448.965 -18.875 ;
        RECT 447.275 -19.205 447.605 -18.875 ;
        RECT 445.915 -19.205 446.245 -18.875 ;
        RECT 444.555 -19.205 444.885 -18.875 ;
        RECT 443.195 -19.205 443.525 -18.875 ;
        RECT 441.835 -19.205 442.165 -18.875 ;
        RECT 440.475 -19.205 440.805 -18.875 ;
        RECT 439.115 -19.205 439.445 -18.875 ;
        RECT 436.395 -19.205 436.725 -18.875 ;
        RECT 433.675 -19.205 434.005 -18.875 ;
        RECT 432.315 -19.205 432.645 -18.875 ;
        RECT 430.955 -19.205 431.285 -18.875 ;
        RECT 429.595 -19.205 429.925 -18.875 ;
        RECT 428.235 -19.205 428.565 -18.875 ;
        RECT 426.875 -19.205 427.205 -18.875 ;
        RECT 425.515 -19.205 425.845 -18.875 ;
        RECT 424.155 -19.205 424.485 -18.875 ;
        RECT 421.435 -19.205 421.765 -18.875 ;
        RECT 418.715 -19.205 419.045 -18.875 ;
        RECT 417.355 -19.205 417.685 -18.875 ;
        RECT 415.995 -19.205 416.325 -18.875 ;
        RECT 414.635 -19.205 414.965 -18.875 ;
        RECT 413.275 -19.205 413.605 -18.875 ;
        RECT 411.915 -19.205 412.245 -18.875 ;
        RECT 410.555 -19.205 410.885 -18.875 ;
        RECT 406.475 -19.205 406.805 -18.875 ;
        RECT 403.755 -19.205 404.085 -18.875 ;
        RECT 402.395 -19.205 402.725 -18.875 ;
        RECT 401.035 -19.205 401.365 -18.875 ;
        RECT 399.675 -19.205 400.005 -18.875 ;
        RECT 398.315 -19.205 398.645 -18.875 ;
        RECT 396.955 -19.205 397.285 -18.875 ;
        RECT 395.595 -19.205 395.925 -18.875 ;
        RECT 391.515 -19.205 391.845 -18.875 ;
        RECT 388.795 -19.205 389.125 -18.875 ;
        RECT 387.435 -19.205 387.765 -18.875 ;
        RECT 386.075 -19.205 386.405 -18.875 ;
        RECT 384.715 -19.205 385.045 -18.875 ;
        RECT 383.355 -19.205 383.685 -18.875 ;
        RECT 381.995 -19.205 382.325 -18.875 ;
        RECT 380.635 -19.205 380.965 -18.875 ;
        RECT 376.555 -19.205 376.885 -18.875 ;
        RECT 373.835 -19.205 374.165 -18.875 ;
        RECT 372.475 -19.205 372.805 -18.875 ;
        RECT 371.115 -19.205 371.445 -18.875 ;
        RECT 369.755 -19.205 370.085 -18.875 ;
        RECT 368.395 -19.205 368.725 -18.875 ;
        RECT 367.035 -19.205 367.365 -18.875 ;
        RECT 365.675 -19.205 366.005 -18.875 ;
        RECT 361.595 -19.205 361.925 -18.875 ;
        RECT 358.875 -19.205 359.205 -18.875 ;
        RECT 357.515 -19.205 357.845 -18.875 ;
        RECT 356.155 -19.205 356.485 -18.875 ;
        RECT 354.795 -19.205 355.125 -18.875 ;
        RECT 353.435 -19.205 353.765 -18.875 ;
        RECT 352.075 -19.205 352.405 -18.875 ;
        RECT 350.715 -19.205 351.045 -18.875 ;
        RECT 346.635 -19.205 346.965 -18.875 ;
        RECT 343.915 -19.205 344.245 -18.875 ;
        RECT 342.555 -19.205 342.885 -18.875 ;
        RECT 341.195 -19.205 341.525 -18.875 ;
        RECT 339.835 -19.205 340.165 -18.875 ;
        RECT 338.475 -19.205 338.805 -18.875 ;
        RECT 337.115 -19.205 337.445 -18.875 ;
        RECT 335.755 -19.205 336.085 -18.875 ;
        RECT 331.675 -19.205 332.005 -18.875 ;
        RECT 328.955 -19.205 329.285 -18.875 ;
        RECT 327.595 -19.205 327.925 -18.875 ;
        RECT 326.235 -19.205 326.565 -18.875 ;
        RECT 324.875 -19.205 325.205 -18.875 ;
        RECT 323.515 -19.205 323.845 -18.875 ;
        RECT 322.155 -19.205 322.485 -18.875 ;
        RECT 320.795 -19.205 321.125 -18.875 ;
        RECT 316.715 -19.205 317.045 -18.875 ;
        RECT 313.995 -19.205 314.325 -18.875 ;
        RECT 312.635 -19.205 312.965 -18.875 ;
        RECT 311.275 -19.205 311.605 -18.875 ;
        RECT 309.915 -19.205 310.245 -18.875 ;
        RECT 308.555 -19.205 308.885 -18.875 ;
        RECT 307.195 -19.205 307.525 -18.875 ;
        RECT 305.835 -19.205 306.165 -18.875 ;
        RECT 300.395 -19.205 300.725 -18.875 ;
        RECT 299.035 -19.205 299.365 -18.875 ;
        RECT 297.675 -19.205 298.005 -18.875 ;
        RECT 296.315 -19.205 296.645 -18.875 ;
        RECT 294.955 -19.205 295.285 -18.875 ;
        RECT 293.595 -19.205 293.925 -18.875 ;
        RECT 292.235 -19.205 292.565 -18.875 ;
        RECT 290.875 -19.205 291.205 -18.875 ;
        RECT 285.435 -19.205 285.765 -18.875 ;
        RECT 284.075 -19.205 284.405 -18.875 ;
        RECT 282.715 -19.205 283.045 -18.875 ;
        RECT 281.355 -19.205 281.685 -18.875 ;
        RECT 279.995 -19.205 280.325 -18.875 ;
        RECT 278.635 -19.205 278.965 -18.875 ;
        RECT 277.275 -19.205 277.605 -18.875 ;
        RECT 275.915 -19.205 276.245 -18.875 ;
        RECT 270.475 -19.205 270.805 -18.875 ;
        RECT 269.115 -19.205 269.445 -18.875 ;
        RECT 267.755 -19.205 268.085 -18.875 ;
        RECT 266.395 -19.205 266.725 -18.875 ;
        RECT 265.035 -19.205 265.365 -18.875 ;
        RECT 263.675 -19.205 264.005 -18.875 ;
        RECT 262.315 -19.205 262.645 -18.875 ;
        RECT 260.955 -19.205 261.285 -18.875 ;
        RECT 255.515 -19.205 255.845 -18.875 ;
        RECT 254.155 -19.205 254.485 -18.875 ;
        RECT 252.795 -19.205 253.125 -18.875 ;
        RECT 251.435 -19.205 251.765 -18.875 ;
        RECT 250.075 -19.205 250.405 -18.875 ;
        RECT 248.715 -19.205 249.045 -18.875 ;
        RECT 247.355 -19.205 247.685 -18.875 ;
        RECT 245.995 -19.205 246.325 -18.875 ;
        RECT 240.555 -19.205 240.885 -18.875 ;
        RECT 239.195 -19.205 239.525 -18.875 ;
        RECT 237.835 -19.205 238.165 -18.875 ;
        RECT 236.475 -19.205 236.805 -18.875 ;
        RECT 235.115 -19.205 235.445 -18.875 ;
        RECT 233.755 -19.205 234.085 -18.875 ;
        RECT 232.395 -19.205 232.725 -18.875 ;
        RECT 231.035 -19.205 231.365 -18.875 ;
        RECT 225.595 -19.205 225.925 -18.875 ;
        RECT 224.235 -19.205 224.565 -18.875 ;
        RECT 222.875 -19.205 223.205 -18.875 ;
        RECT 221.515 -19.205 221.845 -18.875 ;
        RECT 220.155 -19.205 220.485 -18.875 ;
        RECT 218.795 -19.205 219.125 -18.875 ;
        RECT 217.435 -19.205 217.765 -18.875 ;
        RECT 216.075 -19.205 216.405 -18.875 ;
        RECT 210.635 -19.205 210.965 -18.875 ;
        RECT 209.275 -19.205 209.605 -18.875 ;
        RECT 207.915 -19.205 208.245 -18.875 ;
        RECT 206.555 -19.205 206.885 -18.875 ;
        RECT 205.195 -19.205 205.525 -18.875 ;
        RECT 203.835 -19.205 204.165 -18.875 ;
        RECT 202.475 -19.205 202.805 -18.875 ;
        RECT 201.115 -19.205 201.445 -18.875 ;
        RECT 195.675 -19.205 196.005 -18.875 ;
        RECT 194.315 -19.205 194.645 -18.875 ;
        RECT 192.955 -19.205 193.285 -18.875 ;
        RECT 191.595 -19.205 191.925 -18.875 ;
        RECT 190.235 -19.205 190.565 -18.875 ;
        RECT 188.875 -19.205 189.205 -18.875 ;
        RECT 187.515 -19.205 187.845 -18.875 ;
        RECT 186.155 -19.205 186.485 -18.875 ;
        RECT 180.715 -19.205 181.045 -18.875 ;
        RECT 179.355 -19.205 179.685 -18.875 ;
        RECT 177.995 -19.205 178.325 -18.875 ;
        RECT 176.635 -19.205 176.965 -18.875 ;
        RECT 175.275 -19.205 175.605 -18.875 ;
        RECT 173.915 -19.205 174.245 -18.875 ;
        RECT 172.555 -19.205 172.885 -18.875 ;
        RECT 171.195 -19.205 171.525 -18.875 ;
        RECT 165.755 -19.205 166.085 -18.875 ;
        RECT 164.395 -19.205 164.725 -18.875 ;
        RECT 163.035 -19.205 163.365 -18.875 ;
        RECT 161.675 -19.205 162.005 -18.875 ;
        RECT 160.315 -19.205 160.645 -18.875 ;
        RECT 158.955 -19.205 159.285 -18.875 ;
        RECT 157.595 -19.205 157.925 -18.875 ;
        RECT 156.235 -19.205 156.565 -18.875 ;
        RECT 150.795 -19.205 151.125 -18.875 ;
        RECT 149.435 -19.205 149.765 -18.875 ;
        RECT 148.075 -19.205 148.405 -18.875 ;
        RECT 146.715 -19.205 147.045 -18.875 ;
        RECT 145.355 -19.205 145.685 -18.875 ;
        RECT 143.995 -19.205 144.325 -18.875 ;
        RECT 142.635 -19.205 142.965 -18.875 ;
        RECT 141.275 -19.205 141.605 -18.875 ;
        RECT 135.835 -19.205 136.165 -18.875 ;
        RECT 134.475 -19.205 134.805 -18.875 ;
        RECT 133.115 -19.205 133.445 -18.875 ;
        RECT 131.755 -19.205 132.085 -18.875 ;
        RECT 130.395 -19.205 130.725 -18.875 ;
        RECT 129.035 -19.205 129.365 -18.875 ;
        RECT 127.675 -19.205 128.005 -18.875 ;
        RECT 126.315 -19.205 126.645 -18.875 ;
        RECT 120.875 -19.205 121.205 -18.875 ;
        RECT 119.515 -19.205 119.845 -18.875 ;
        RECT 118.155 -19.205 118.485 -18.875 ;
        RECT 116.795 -19.205 117.125 -18.875 ;
        RECT 115.435 -19.205 115.765 -18.875 ;
        RECT 114.075 -19.205 114.405 -18.875 ;
        RECT 112.715 -19.205 113.045 -18.875 ;
        RECT 111.355 -19.205 111.685 -18.875 ;
        RECT 105.915 -19.205 106.245 -18.875 ;
        RECT 104.555 -19.205 104.885 -18.875 ;
        RECT 103.195 -19.205 103.525 -18.875 ;
        RECT 101.835 -19.205 102.165 -18.875 ;
        RECT 100.475 -19.205 100.805 -18.875 ;
        RECT 99.115 -19.205 99.445 -18.875 ;
        RECT 97.755 -19.205 98.085 -18.875 ;
        RECT 96.395 -19.205 96.725 -18.875 ;
        RECT 93.675 -19.205 94.005 -18.875 ;
        RECT 90.955 -19.205 91.285 -18.875 ;
        RECT 89.595 -19.205 89.925 -18.875 ;
        RECT 88.235 -19.205 88.565 -18.875 ;
        RECT 86.875 -19.205 87.205 -18.875 ;
        RECT 85.515 -19.205 85.845 -18.875 ;
        RECT 84.155 -19.205 84.485 -18.875 ;
        RECT 82.795 -19.205 83.125 -18.875 ;
        RECT 81.435 -19.205 81.765 -18.875 ;
        RECT 78.715 -19.205 79.045 -18.875 ;
        RECT 75.995 -19.205 76.325 -18.875 ;
        RECT 74.635 -19.205 74.965 -18.875 ;
        RECT 73.275 -19.205 73.605 -18.875 ;
        RECT 71.915 -19.205 72.245 -18.875 ;
        RECT 70.555 -19.205 70.885 -18.875 ;
        RECT 69.195 -19.205 69.525 -18.875 ;
        RECT 67.835 -19.205 68.165 -18.875 ;
        RECT 63.755 -19.205 64.085 -18.875 ;
        RECT 61.035 -19.205 61.365 -18.875 ;
        RECT 59.675 -19.205 60.005 -18.875 ;
        RECT 58.315 -19.205 58.645 -18.875 ;
        RECT 56.955 -19.205 57.285 -18.875 ;
        RECT 55.595 -19.205 55.925 -18.875 ;
        RECT 54.235 -19.205 54.565 -18.875 ;
        RECT 52.875 -19.205 53.205 -18.875 ;
        RECT 48.795 -19.205 49.125 -18.875 ;
        RECT 46.075 -19.205 46.405 -18.875 ;
        RECT 44.715 -19.205 45.045 -18.875 ;
        RECT 43.355 -19.205 43.685 -18.875 ;
        RECT 41.995 -19.205 42.325 -18.875 ;
        RECT 40.635 -19.205 40.965 -18.875 ;
        RECT 39.275 -19.205 39.605 -18.875 ;
        RECT 37.915 -19.205 38.245 -18.875 ;
        RECT 33.835 -19.205 34.165 -18.875 ;
        RECT 31.115 -19.205 31.445 -18.875 ;
        RECT 29.755 -19.205 30.085 -18.875 ;
        RECT 28.395 -19.205 28.725 -18.875 ;
        RECT 27.035 -19.205 27.365 -18.875 ;
        RECT 25.675 -19.205 26.005 -18.875 ;
        RECT 24.315 -19.205 24.645 -18.875 ;
        RECT 22.955 -19.205 23.285 -18.875 ;
        RECT 18.875 -19.205 19.205 -18.875 ;
        RECT 16.155 -19.205 16.485 -18.875 ;
        RECT 14.795 -19.205 15.125 -18.875 ;
        RECT 13.435 -19.205 13.765 -18.875 ;
        RECT 12.075 -19.205 12.405 -18.875 ;
        RECT 954.555 -19.205 954.885 -18.875 ;
        RECT 920.555 -19.2 954.885 -18.88 ;
        RECT 953.195 -19.205 953.525 -18.875 ;
        RECT 951.835 -19.205 952.165 -18.875 ;
        RECT 950.475 -19.205 950.805 -18.875 ;
        RECT 949.115 -19.205 949.445 -18.875 ;
        RECT 947.755 -19.205 948.085 -18.875 ;
        RECT 946.395 -19.205 946.725 -18.875 ;
        RECT 945.035 -19.205 945.365 -18.875 ;
        RECT 940.955 -19.205 941.285 -18.875 ;
        RECT 939.595 -19.205 939.925 -18.875 ;
        RECT 938.235 -19.205 938.565 -18.875 ;
        RECT 936.875 -19.205 937.205 -18.875 ;
        RECT 935.515 -19.205 935.845 -18.875 ;
        RECT 934.155 -19.205 934.485 -18.875 ;
        RECT 932.795 -19.205 933.125 -18.875 ;
        RECT 931.435 -19.205 931.765 -18.875 ;
        RECT 925.995 -19.205 926.325 -18.875 ;
        RECT 924.635 -19.205 924.965 -18.875 ;
        RECT 923.275 -19.205 923.605 -18.875 ;
        RECT 921.915 -19.205 922.245 -18.875 ;
        RECT 920.555 -19.205 920.885 -18.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -15.12 678.475 -14.8 ;
        RECT 677.115 -15.125 677.445 -14.795 ;
        RECT 675.755 -15.125 676.085 -14.795 ;
        RECT 674.395 -15.125 674.725 -14.795 ;
        RECT 673.035 -15.125 673.365 -14.795 ;
        RECT 671.675 -15.125 672.005 -14.795 ;
        RECT 670.315 -15.125 670.645 -14.795 ;
        RECT 668.955 -15.125 669.285 -14.795 ;
        RECT 667.595 -15.125 667.925 -14.795 ;
        RECT 666.235 -15.125 666.565 -14.795 ;
        RECT 664.875 -15.125 665.205 -14.795 ;
        RECT 663.515 -15.125 663.845 -14.795 ;
        RECT 662.155 -15.125 662.485 -14.795 ;
        RECT 660.795 -15.125 661.125 -14.795 ;
        RECT 659.435 -15.125 659.765 -14.795 ;
        RECT 658.075 -15.125 658.405 -14.795 ;
        RECT 656.715 -15.125 657.045 -14.795 ;
        RECT 655.355 -15.125 655.685 -14.795 ;
        RECT 653.995 -15.125 654.325 -14.795 ;
        RECT 652.635 -15.125 652.965 -14.795 ;
        RECT 651.275 -15.125 651.605 -14.795 ;
        RECT 649.915 -15.125 650.245 -14.795 ;
        RECT 648.555 -15.125 648.885 -14.795 ;
        RECT 647.195 -15.125 647.525 -14.795 ;
        RECT 645.835 -15.125 646.165 -14.795 ;
        RECT 644.475 -15.125 644.805 -14.795 ;
        RECT 643.115 -15.125 643.445 -14.795 ;
        RECT 641.755 -15.125 642.085 -14.795 ;
        RECT 640.395 -15.125 640.725 -14.795 ;
        RECT 639.035 -15.125 639.365 -14.795 ;
        RECT 637.675 -15.125 638.005 -14.795 ;
        RECT 636.315 -15.125 636.645 -14.795 ;
        RECT 634.955 -15.125 635.285 -14.795 ;
        RECT 633.595 -15.125 633.925 -14.795 ;
        RECT 632.235 -15.125 632.565 -14.795 ;
        RECT 630.875 -15.125 631.205 -14.795 ;
        RECT 629.515 -15.125 629.845 -14.795 ;
        RECT 628.155 -15.125 628.485 -14.795 ;
        RECT 626.795 -15.125 627.125 -14.795 ;
        RECT 625.435 -15.125 625.765 -14.795 ;
        RECT 624.075 -15.125 624.405 -14.795 ;
        RECT 622.715 -15.125 623.045 -14.795 ;
        RECT 621.355 -15.125 621.685 -14.795 ;
        RECT 619.995 -15.125 620.325 -14.795 ;
        RECT 618.635 -15.125 618.965 -14.795 ;
        RECT 617.275 -15.125 617.605 -14.795 ;
        RECT 615.915 -15.125 616.245 -14.795 ;
        RECT 614.555 -15.125 614.885 -14.795 ;
        RECT 613.195 -15.125 613.525 -14.795 ;
        RECT 611.835 -15.125 612.165 -14.795 ;
        RECT 610.475 -15.125 610.805 -14.795 ;
        RECT 609.115 -15.125 609.445 -14.795 ;
        RECT 607.755 -15.125 608.085 -14.795 ;
        RECT 606.395 -15.125 606.725 -14.795 ;
        RECT 605.035 -15.125 605.365 -14.795 ;
        RECT 603.675 -15.125 604.005 -14.795 ;
        RECT 602.315 -15.125 602.645 -14.795 ;
        RECT 600.955 -15.125 601.285 -14.795 ;
        RECT 599.595 -15.125 599.925 -14.795 ;
        RECT 598.235 -15.125 598.565 -14.795 ;
        RECT 596.875 -15.125 597.205 -14.795 ;
        RECT 595.515 -15.125 595.845 -14.795 ;
        RECT 594.155 -15.125 594.485 -14.795 ;
        RECT 592.795 -15.125 593.125 -14.795 ;
        RECT 591.435 -15.125 591.765 -14.795 ;
        RECT 590.075 -15.125 590.405 -14.795 ;
        RECT 588.715 -15.125 589.045 -14.795 ;
        RECT 587.355 -15.125 587.685 -14.795 ;
        RECT 585.995 -15.125 586.325 -14.795 ;
        RECT 584.635 -15.125 584.965 -14.795 ;
        RECT 583.275 -15.125 583.605 -14.795 ;
        RECT 581.915 -15.125 582.245 -14.795 ;
        RECT 580.555 -15.125 580.885 -14.795 ;
        RECT 579.195 -15.125 579.525 -14.795 ;
        RECT 577.835 -15.125 578.165 -14.795 ;
        RECT 576.475 -15.125 576.805 -14.795 ;
        RECT 575.115 -15.125 575.445 -14.795 ;
        RECT 573.755 -15.125 574.085 -14.795 ;
        RECT 572.395 -15.125 572.725 -14.795 ;
        RECT 571.035 -15.125 571.365 -14.795 ;
        RECT 569.675 -15.125 570.005 -14.795 ;
        RECT 568.315 -15.125 568.645 -14.795 ;
        RECT 566.955 -15.125 567.285 -14.795 ;
        RECT 565.595 -15.125 565.925 -14.795 ;
        RECT 564.235 -15.125 564.565 -14.795 ;
        RECT 562.875 -15.125 563.205 -14.795 ;
        RECT 561.515 -15.125 561.845 -14.795 ;
        RECT 560.155 -15.125 560.485 -14.795 ;
        RECT 558.795 -15.125 559.125 -14.795 ;
        RECT 557.435 -15.125 557.765 -14.795 ;
        RECT 556.075 -15.125 556.405 -14.795 ;
        RECT 554.715 -15.125 555.045 -14.795 ;
        RECT 553.355 -15.125 553.685 -14.795 ;
        RECT 551.995 -15.125 552.325 -14.795 ;
        RECT 550.635 -15.125 550.965 -14.795 ;
        RECT 549.275 -15.125 549.605 -14.795 ;
        RECT 547.915 -15.125 548.245 -14.795 ;
        RECT 546.555 -15.125 546.885 -14.795 ;
        RECT 545.195 -15.125 545.525 -14.795 ;
        RECT 543.835 -15.125 544.165 -14.795 ;
        RECT 542.475 -15.125 542.805 -14.795 ;
        RECT 541.115 -15.125 541.445 -14.795 ;
        RECT 539.755 -15.125 540.085 -14.795 ;
        RECT 538.395 -15.125 538.725 -14.795 ;
        RECT 537.035 -15.125 537.365 -14.795 ;
        RECT 535.675 -15.125 536.005 -14.795 ;
        RECT 534.315 -15.125 534.645 -14.795 ;
        RECT 532.955 -15.125 533.285 -14.795 ;
        RECT 531.595 -15.125 531.925 -14.795 ;
        RECT 530.235 -15.125 530.565 -14.795 ;
        RECT 528.875 -15.125 529.205 -14.795 ;
        RECT 527.515 -15.125 527.845 -14.795 ;
        RECT 526.155 -15.125 526.485 -14.795 ;
        RECT 524.795 -15.125 525.125 -14.795 ;
        RECT 523.435 -15.125 523.765 -14.795 ;
        RECT 522.075 -15.125 522.405 -14.795 ;
        RECT 520.715 -15.125 521.045 -14.795 ;
        RECT 519.355 -15.125 519.685 -14.795 ;
        RECT 517.995 -15.125 518.325 -14.795 ;
        RECT 516.635 -15.125 516.965 -14.795 ;
        RECT 515.275 -15.125 515.605 -14.795 ;
        RECT 513.915 -15.125 514.245 -14.795 ;
        RECT 512.555 -15.125 512.885 -14.795 ;
        RECT 511.195 -15.125 511.525 -14.795 ;
        RECT 509.835 -15.125 510.165 -14.795 ;
        RECT 508.475 -15.125 508.805 -14.795 ;
        RECT 507.115 -15.125 507.445 -14.795 ;
        RECT 505.755 -15.125 506.085 -14.795 ;
        RECT 504.395 -15.125 504.725 -14.795 ;
        RECT 503.035 -15.125 503.365 -14.795 ;
        RECT 501.675 -15.125 502.005 -14.795 ;
        RECT 500.315 -15.125 500.645 -14.795 ;
        RECT 498.955 -15.125 499.285 -14.795 ;
        RECT 497.595 -15.125 497.925 -14.795 ;
        RECT 496.235 -15.125 496.565 -14.795 ;
        RECT 494.875 -15.125 495.205 -14.795 ;
        RECT 493.515 -15.125 493.845 -14.795 ;
        RECT 492.155 -15.125 492.485 -14.795 ;
        RECT 490.795 -15.125 491.125 -14.795 ;
        RECT 489.435 -15.125 489.765 -14.795 ;
        RECT 488.075 -15.125 488.405 -14.795 ;
        RECT 486.715 -15.125 487.045 -14.795 ;
        RECT 485.355 -15.125 485.685 -14.795 ;
        RECT 483.995 -15.125 484.325 -14.795 ;
        RECT 482.635 -15.125 482.965 -14.795 ;
        RECT 481.275 -15.125 481.605 -14.795 ;
        RECT 479.915 -15.125 480.245 -14.795 ;
        RECT 478.555 -15.125 478.885 -14.795 ;
        RECT 477.195 -15.125 477.525 -14.795 ;
        RECT 475.835 -15.125 476.165 -14.795 ;
        RECT 474.475 -15.125 474.805 -14.795 ;
        RECT 473.115 -15.125 473.445 -14.795 ;
        RECT 471.755 -15.125 472.085 -14.795 ;
        RECT 470.395 -15.125 470.725 -14.795 ;
        RECT 469.035 -15.125 469.365 -14.795 ;
        RECT 467.675 -15.125 468.005 -14.795 ;
        RECT 466.315 -15.125 466.645 -14.795 ;
        RECT 464.955 -15.125 465.285 -14.795 ;
        RECT 463.595 -15.125 463.925 -14.795 ;
        RECT 462.235 -15.125 462.565 -14.795 ;
        RECT 460.875 -15.125 461.205 -14.795 ;
        RECT 459.515 -15.125 459.845 -14.795 ;
        RECT 458.155 -15.125 458.485 -14.795 ;
        RECT 456.795 -15.125 457.125 -14.795 ;
        RECT 455.435 -15.125 455.765 -14.795 ;
        RECT 454.075 -15.125 454.405 -14.795 ;
        RECT 452.715 -15.125 453.045 -14.795 ;
        RECT 451.355 -15.125 451.685 -14.795 ;
        RECT 449.995 -15.125 450.325 -14.795 ;
        RECT 448.635 -15.125 448.965 -14.795 ;
        RECT 447.275 -15.125 447.605 -14.795 ;
        RECT 445.915 -15.125 446.245 -14.795 ;
        RECT 444.555 -15.125 444.885 -14.795 ;
        RECT 443.195 -15.125 443.525 -14.795 ;
        RECT 441.835 -15.125 442.165 -14.795 ;
        RECT 440.475 -15.125 440.805 -14.795 ;
        RECT 439.115 -15.125 439.445 -14.795 ;
        RECT 437.755 -15.125 438.085 -14.795 ;
        RECT 436.395 -15.125 436.725 -14.795 ;
        RECT 435.035 -15.125 435.365 -14.795 ;
        RECT 433.675 -15.125 434.005 -14.795 ;
        RECT 432.315 -15.125 432.645 -14.795 ;
        RECT 430.955 -15.125 431.285 -14.795 ;
        RECT 429.595 -15.125 429.925 -14.795 ;
        RECT 428.235 -15.125 428.565 -14.795 ;
        RECT 426.875 -15.125 427.205 -14.795 ;
        RECT 425.515 -15.125 425.845 -14.795 ;
        RECT 424.155 -15.125 424.485 -14.795 ;
        RECT 422.795 -15.125 423.125 -14.795 ;
        RECT 421.435 -15.125 421.765 -14.795 ;
        RECT 420.075 -15.125 420.405 -14.795 ;
        RECT 418.715 -15.125 419.045 -14.795 ;
        RECT 417.355 -15.125 417.685 -14.795 ;
        RECT 415.995 -15.125 416.325 -14.795 ;
        RECT 414.635 -15.125 414.965 -14.795 ;
        RECT 413.275 -15.125 413.605 -14.795 ;
        RECT 411.915 -15.125 412.245 -14.795 ;
        RECT 410.555 -15.125 410.885 -14.795 ;
        RECT 409.195 -15.125 409.525 -14.795 ;
        RECT 407.835 -15.125 408.165 -14.795 ;
        RECT 406.475 -15.125 406.805 -14.795 ;
        RECT 405.115 -15.125 405.445 -14.795 ;
        RECT 403.755 -15.125 404.085 -14.795 ;
        RECT 402.395 -15.125 402.725 -14.795 ;
        RECT 401.035 -15.125 401.365 -14.795 ;
        RECT 399.675 -15.125 400.005 -14.795 ;
        RECT 398.315 -15.125 398.645 -14.795 ;
        RECT 396.955 -15.125 397.285 -14.795 ;
        RECT 395.595 -15.125 395.925 -14.795 ;
        RECT 394.235 -15.125 394.565 -14.795 ;
        RECT 392.875 -15.125 393.205 -14.795 ;
        RECT 391.515 -15.125 391.845 -14.795 ;
        RECT 390.155 -15.125 390.485 -14.795 ;
        RECT 388.795 -15.125 389.125 -14.795 ;
        RECT 387.435 -15.125 387.765 -14.795 ;
        RECT 386.075 -15.125 386.405 -14.795 ;
        RECT 384.715 -15.125 385.045 -14.795 ;
        RECT 383.355 -15.125 383.685 -14.795 ;
        RECT 381.995 -15.125 382.325 -14.795 ;
        RECT 380.635 -15.125 380.965 -14.795 ;
        RECT 379.275 -15.125 379.605 -14.795 ;
        RECT 377.915 -15.125 378.245 -14.795 ;
        RECT 376.555 -15.125 376.885 -14.795 ;
        RECT 375.195 -15.125 375.525 -14.795 ;
        RECT 373.835 -15.125 374.165 -14.795 ;
        RECT 372.475 -15.125 372.805 -14.795 ;
        RECT 371.115 -15.125 371.445 -14.795 ;
        RECT 369.755 -15.125 370.085 -14.795 ;
        RECT 368.395 -15.125 368.725 -14.795 ;
        RECT 367.035 -15.125 367.365 -14.795 ;
        RECT 365.675 -15.125 366.005 -14.795 ;
        RECT 364.315 -15.125 364.645 -14.795 ;
        RECT 362.955 -15.125 363.285 -14.795 ;
        RECT 361.595 -15.125 361.925 -14.795 ;
        RECT 360.235 -15.125 360.565 -14.795 ;
        RECT 358.875 -15.125 359.205 -14.795 ;
        RECT 357.515 -15.125 357.845 -14.795 ;
        RECT 356.155 -15.125 356.485 -14.795 ;
        RECT 354.795 -15.125 355.125 -14.795 ;
        RECT 353.435 -15.125 353.765 -14.795 ;
        RECT 352.075 -15.125 352.405 -14.795 ;
        RECT 350.715 -15.125 351.045 -14.795 ;
        RECT 349.355 -15.125 349.685 -14.795 ;
        RECT 347.995 -15.125 348.325 -14.795 ;
        RECT 346.635 -15.125 346.965 -14.795 ;
        RECT 345.275 -15.125 345.605 -14.795 ;
        RECT 343.915 -15.125 344.245 -14.795 ;
        RECT 342.555 -15.125 342.885 -14.795 ;
        RECT 341.195 -15.125 341.525 -14.795 ;
        RECT 339.835 -15.125 340.165 -14.795 ;
        RECT 338.475 -15.125 338.805 -14.795 ;
        RECT 337.115 -15.125 337.445 -14.795 ;
        RECT 335.755 -15.125 336.085 -14.795 ;
        RECT 334.395 -15.125 334.725 -14.795 ;
        RECT 333.035 -15.125 333.365 -14.795 ;
        RECT 331.675 -15.125 332.005 -14.795 ;
        RECT 330.315 -15.125 330.645 -14.795 ;
        RECT 328.955 -15.125 329.285 -14.795 ;
        RECT 327.595 -15.125 327.925 -14.795 ;
        RECT 326.235 -15.125 326.565 -14.795 ;
        RECT 324.875 -15.125 325.205 -14.795 ;
        RECT 323.515 -15.125 323.845 -14.795 ;
        RECT 322.155 -15.125 322.485 -14.795 ;
        RECT 320.795 -15.125 321.125 -14.795 ;
        RECT 319.435 -15.125 319.765 -14.795 ;
        RECT 318.075 -15.125 318.405 -14.795 ;
        RECT 316.715 -15.125 317.045 -14.795 ;
        RECT 315.355 -15.125 315.685 -14.795 ;
        RECT 313.995 -15.125 314.325 -14.795 ;
        RECT 312.635 -15.125 312.965 -14.795 ;
        RECT 311.275 -15.125 311.605 -14.795 ;
        RECT 309.915 -15.125 310.245 -14.795 ;
        RECT 308.555 -15.125 308.885 -14.795 ;
        RECT 307.195 -15.125 307.525 -14.795 ;
        RECT 305.835 -15.125 306.165 -14.795 ;
        RECT 304.475 -15.125 304.805 -14.795 ;
        RECT 303.115 -15.125 303.445 -14.795 ;
        RECT 301.755 -15.125 302.085 -14.795 ;
        RECT 300.395 -15.125 300.725 -14.795 ;
        RECT 299.035 -15.125 299.365 -14.795 ;
        RECT 297.675 -15.125 298.005 -14.795 ;
        RECT 296.315 -15.125 296.645 -14.795 ;
        RECT 294.955 -15.125 295.285 -14.795 ;
        RECT 293.595 -15.125 293.925 -14.795 ;
        RECT 292.235 -15.125 292.565 -14.795 ;
        RECT 290.875 -15.125 291.205 -14.795 ;
        RECT 289.515 -15.125 289.845 -14.795 ;
        RECT 288.155 -15.125 288.485 -14.795 ;
        RECT 286.795 -15.125 287.125 -14.795 ;
        RECT 285.435 -15.125 285.765 -14.795 ;
        RECT 284.075 -15.125 284.405 -14.795 ;
        RECT 282.715 -15.125 283.045 -14.795 ;
        RECT 281.355 -15.125 281.685 -14.795 ;
        RECT 279.995 -15.125 280.325 -14.795 ;
        RECT 278.635 -15.125 278.965 -14.795 ;
        RECT 277.275 -15.125 277.605 -14.795 ;
        RECT 275.915 -15.125 276.245 -14.795 ;
        RECT 274.555 -15.125 274.885 -14.795 ;
        RECT 273.195 -15.125 273.525 -14.795 ;
        RECT 271.835 -15.125 272.165 -14.795 ;
        RECT 270.475 -15.125 270.805 -14.795 ;
        RECT 269.115 -15.125 269.445 -14.795 ;
        RECT 267.755 -15.125 268.085 -14.795 ;
        RECT 266.395 -15.125 266.725 -14.795 ;
        RECT 265.035 -15.125 265.365 -14.795 ;
        RECT 263.675 -15.125 264.005 -14.795 ;
        RECT 262.315 -15.125 262.645 -14.795 ;
        RECT 260.955 -15.125 261.285 -14.795 ;
        RECT 259.595 -15.125 259.925 -14.795 ;
        RECT 258.235 -15.125 258.565 -14.795 ;
        RECT 256.875 -15.125 257.205 -14.795 ;
        RECT 255.515 -15.125 255.845 -14.795 ;
        RECT 254.155 -15.125 254.485 -14.795 ;
        RECT 252.795 -15.125 253.125 -14.795 ;
        RECT 251.435 -15.125 251.765 -14.795 ;
        RECT 250.075 -15.125 250.405 -14.795 ;
        RECT 248.715 -15.125 249.045 -14.795 ;
        RECT 247.355 -15.125 247.685 -14.795 ;
        RECT 245.995 -15.125 246.325 -14.795 ;
        RECT 244.635 -15.125 244.965 -14.795 ;
        RECT 243.275 -15.125 243.605 -14.795 ;
        RECT 241.915 -15.125 242.245 -14.795 ;
        RECT 240.555 -15.125 240.885 -14.795 ;
        RECT 239.195 -15.125 239.525 -14.795 ;
        RECT 237.835 -15.125 238.165 -14.795 ;
        RECT 236.475 -15.125 236.805 -14.795 ;
        RECT 235.115 -15.125 235.445 -14.795 ;
        RECT 233.755 -15.125 234.085 -14.795 ;
        RECT 232.395 -15.125 232.725 -14.795 ;
        RECT 231.035 -15.125 231.365 -14.795 ;
        RECT 229.675 -15.125 230.005 -14.795 ;
        RECT 228.315 -15.125 228.645 -14.795 ;
        RECT 226.955 -15.125 227.285 -14.795 ;
        RECT 225.595 -15.125 225.925 -14.795 ;
        RECT 224.235 -15.125 224.565 -14.795 ;
        RECT 222.875 -15.125 223.205 -14.795 ;
        RECT 221.515 -15.125 221.845 -14.795 ;
        RECT 220.155 -15.125 220.485 -14.795 ;
        RECT 218.795 -15.125 219.125 -14.795 ;
        RECT 217.435 -15.125 217.765 -14.795 ;
        RECT 216.075 -15.125 216.405 -14.795 ;
        RECT 214.715 -15.125 215.045 -14.795 ;
        RECT 213.355 -15.125 213.685 -14.795 ;
        RECT 211.995 -15.125 212.325 -14.795 ;
        RECT 210.635 -15.125 210.965 -14.795 ;
        RECT 209.275 -15.125 209.605 -14.795 ;
        RECT 207.915 -15.125 208.245 -14.795 ;
        RECT 206.555 -15.125 206.885 -14.795 ;
        RECT 205.195 -15.125 205.525 -14.795 ;
        RECT 203.835 -15.125 204.165 -14.795 ;
        RECT 202.475 -15.125 202.805 -14.795 ;
        RECT 201.115 -15.125 201.445 -14.795 ;
        RECT 199.755 -15.125 200.085 -14.795 ;
        RECT 198.395 -15.125 198.725 -14.795 ;
        RECT 197.035 -15.125 197.365 -14.795 ;
        RECT 195.675 -15.125 196.005 -14.795 ;
        RECT 194.315 -15.125 194.645 -14.795 ;
        RECT 192.955 -15.125 193.285 -14.795 ;
        RECT 191.595 -15.125 191.925 -14.795 ;
        RECT 190.235 -15.125 190.565 -14.795 ;
        RECT 188.875 -15.125 189.205 -14.795 ;
        RECT 187.515 -15.125 187.845 -14.795 ;
        RECT 186.155 -15.125 186.485 -14.795 ;
        RECT 184.795 -15.125 185.125 -14.795 ;
        RECT 183.435 -15.125 183.765 -14.795 ;
        RECT 182.075 -15.125 182.405 -14.795 ;
        RECT 180.715 -15.125 181.045 -14.795 ;
        RECT 179.355 -15.125 179.685 -14.795 ;
        RECT 177.995 -15.125 178.325 -14.795 ;
        RECT 176.635 -15.125 176.965 -14.795 ;
        RECT 175.275 -15.125 175.605 -14.795 ;
        RECT 173.915 -15.125 174.245 -14.795 ;
        RECT 172.555 -15.125 172.885 -14.795 ;
        RECT 171.195 -15.125 171.525 -14.795 ;
        RECT 169.835 -15.125 170.165 -14.795 ;
        RECT 168.475 -15.125 168.805 -14.795 ;
        RECT 167.115 -15.125 167.445 -14.795 ;
        RECT 165.755 -15.125 166.085 -14.795 ;
        RECT 164.395 -15.125 164.725 -14.795 ;
        RECT 163.035 -15.125 163.365 -14.795 ;
        RECT 161.675 -15.125 162.005 -14.795 ;
        RECT 160.315 -15.125 160.645 -14.795 ;
        RECT 158.955 -15.125 159.285 -14.795 ;
        RECT 157.595 -15.125 157.925 -14.795 ;
        RECT 156.235 -15.125 156.565 -14.795 ;
        RECT 154.875 -15.125 155.205 -14.795 ;
        RECT 153.515 -15.125 153.845 -14.795 ;
        RECT 152.155 -15.125 152.485 -14.795 ;
        RECT 150.795 -15.125 151.125 -14.795 ;
        RECT 149.435 -15.125 149.765 -14.795 ;
        RECT 148.075 -15.125 148.405 -14.795 ;
        RECT 146.715 -15.125 147.045 -14.795 ;
        RECT 145.355 -15.125 145.685 -14.795 ;
        RECT 143.995 -15.125 144.325 -14.795 ;
        RECT 142.635 -15.125 142.965 -14.795 ;
        RECT 141.275 -15.125 141.605 -14.795 ;
        RECT 139.915 -15.125 140.245 -14.795 ;
        RECT 138.555 -15.125 138.885 -14.795 ;
        RECT 137.195 -15.125 137.525 -14.795 ;
        RECT 135.835 -15.125 136.165 -14.795 ;
        RECT 134.475 -15.125 134.805 -14.795 ;
        RECT 133.115 -15.125 133.445 -14.795 ;
        RECT 131.755 -15.125 132.085 -14.795 ;
        RECT 130.395 -15.125 130.725 -14.795 ;
        RECT 129.035 -15.125 129.365 -14.795 ;
        RECT 127.675 -15.125 128.005 -14.795 ;
        RECT 126.315 -15.125 126.645 -14.795 ;
        RECT 124.955 -15.125 125.285 -14.795 ;
        RECT 123.595 -15.125 123.925 -14.795 ;
        RECT 122.235 -15.125 122.565 -14.795 ;
        RECT 120.875 -15.125 121.205 -14.795 ;
        RECT 119.515 -15.125 119.845 -14.795 ;
        RECT 118.155 -15.125 118.485 -14.795 ;
        RECT 116.795 -15.125 117.125 -14.795 ;
        RECT 115.435 -15.125 115.765 -14.795 ;
        RECT 114.075 -15.125 114.405 -14.795 ;
        RECT 112.715 -15.125 113.045 -14.795 ;
        RECT 111.355 -15.125 111.685 -14.795 ;
        RECT 109.995 -15.125 110.325 -14.795 ;
        RECT 108.635 -15.125 108.965 -14.795 ;
        RECT 107.275 -15.125 107.605 -14.795 ;
        RECT 105.915 -15.125 106.245 -14.795 ;
        RECT 104.555 -15.125 104.885 -14.795 ;
        RECT 103.195 -15.125 103.525 -14.795 ;
        RECT 101.835 -15.125 102.165 -14.795 ;
        RECT 100.475 -15.125 100.805 -14.795 ;
        RECT 99.115 -15.125 99.445 -14.795 ;
        RECT 97.755 -15.125 98.085 -14.795 ;
        RECT 96.395 -15.125 96.725 -14.795 ;
        RECT 95.035 -15.125 95.365 -14.795 ;
        RECT 93.675 -15.125 94.005 -14.795 ;
        RECT 92.315 -15.125 92.645 -14.795 ;
        RECT 90.955 -15.125 91.285 -14.795 ;
        RECT 89.595 -15.125 89.925 -14.795 ;
        RECT 88.235 -15.125 88.565 -14.795 ;
        RECT 86.875 -15.125 87.205 -14.795 ;
        RECT 85.515 -15.125 85.845 -14.795 ;
        RECT 84.155 -15.125 84.485 -14.795 ;
        RECT 82.795 -15.125 83.125 -14.795 ;
        RECT 81.435 -15.125 81.765 -14.795 ;
        RECT 80.075 -15.125 80.405 -14.795 ;
        RECT 78.715 -15.125 79.045 -14.795 ;
        RECT 77.355 -15.125 77.685 -14.795 ;
        RECT 75.995 -15.125 76.325 -14.795 ;
        RECT 74.635 -15.125 74.965 -14.795 ;
        RECT 73.275 -15.125 73.605 -14.795 ;
        RECT 71.915 -15.125 72.245 -14.795 ;
        RECT 70.555 -15.125 70.885 -14.795 ;
        RECT 69.195 -15.125 69.525 -14.795 ;
        RECT 67.835 -15.125 68.165 -14.795 ;
        RECT 66.475 -15.125 66.805 -14.795 ;
        RECT 65.115 -15.125 65.445 -14.795 ;
        RECT 63.755 -15.125 64.085 -14.795 ;
        RECT 62.395 -15.125 62.725 -14.795 ;
        RECT 61.035 -15.125 61.365 -14.795 ;
        RECT 59.675 -15.125 60.005 -14.795 ;
        RECT 58.315 -15.125 58.645 -14.795 ;
        RECT 56.955 -15.125 57.285 -14.795 ;
        RECT 55.595 -15.125 55.925 -14.795 ;
        RECT 54.235 -15.125 54.565 -14.795 ;
        RECT 52.875 -15.125 53.205 -14.795 ;
        RECT 51.515 -15.125 51.845 -14.795 ;
        RECT 50.155 -15.125 50.485 -14.795 ;
        RECT 48.795 -15.125 49.125 -14.795 ;
        RECT 47.435 -15.125 47.765 -14.795 ;
        RECT 46.075 -15.125 46.405 -14.795 ;
        RECT 44.715 -15.125 45.045 -14.795 ;
        RECT 43.355 -15.125 43.685 -14.795 ;
        RECT 41.995 -15.125 42.325 -14.795 ;
        RECT 40.635 -15.125 40.965 -14.795 ;
        RECT 39.275 -15.125 39.605 -14.795 ;
        RECT 37.915 -15.125 38.245 -14.795 ;
        RECT 36.555 -15.125 36.885 -14.795 ;
        RECT 35.195 -15.125 35.525 -14.795 ;
        RECT 33.835 -15.125 34.165 -14.795 ;
        RECT 32.475 -15.125 32.805 -14.795 ;
        RECT 31.115 -15.125 31.445 -14.795 ;
        RECT 29.755 -15.125 30.085 -14.795 ;
        RECT 28.395 -15.125 28.725 -14.795 ;
        RECT 27.035 -15.125 27.365 -14.795 ;
        RECT 25.675 -15.125 26.005 -14.795 ;
        RECT 24.315 -15.125 24.645 -14.795 ;
        RECT 22.955 -15.125 23.285 -14.795 ;
        RECT 21.595 -15.125 21.925 -14.795 ;
        RECT 20.235 -15.125 20.565 -14.795 ;
        RECT 18.875 -15.125 19.205 -14.795 ;
        RECT 17.515 -15.125 17.845 -14.795 ;
        RECT 16.155 -15.125 16.485 -14.795 ;
        RECT 14.795 -15.125 15.125 -14.795 ;
        RECT 13.435 -15.125 13.765 -14.795 ;
        RECT 12.075 -15.125 12.405 -14.795 ;
        RECT 10.715 -15.125 11.045 -14.795 ;
        RECT 9.355 -15.125 9.685 -14.795 ;
        RECT 7.995 -15.125 8.325 -14.795 ;
        RECT 6.635 -15.125 6.965 -14.795 ;
        RECT 5.275 -15.125 5.605 -14.795 ;
        RECT 3.915 -15.125 4.245 -14.795 ;
        RECT 2.555 -15.125 2.885 -14.795 ;
        RECT 1.195 -15.125 1.525 -14.795 ;
        RECT -0.165 -15.125 0.165 -14.795 ;
        RECT -1.525 -15.125 -1.195 -14.795 ;
        RECT 954.555 -15.125 954.885 -14.795 ;
        RECT 678.475 -15.12 954.885 -14.8 ;
        RECT 953.195 -15.125 953.525 -14.795 ;
        RECT 951.835 -15.125 952.165 -14.795 ;
        RECT 950.475 -15.125 950.805 -14.795 ;
        RECT 949.115 -15.125 949.445 -14.795 ;
        RECT 947.755 -15.125 948.085 -14.795 ;
        RECT 946.395 -15.125 946.725 -14.795 ;
        RECT 945.035 -15.125 945.365 -14.795 ;
        RECT 943.675 -15.125 944.005 -14.795 ;
        RECT 942.315 -15.125 942.645 -14.795 ;
        RECT 940.955 -15.125 941.285 -14.795 ;
        RECT 939.595 -15.125 939.925 -14.795 ;
        RECT 938.235 -15.125 938.565 -14.795 ;
        RECT 936.875 -15.125 937.205 -14.795 ;
        RECT 935.515 -15.125 935.845 -14.795 ;
        RECT 934.155 -15.125 934.485 -14.795 ;
        RECT 932.795 -15.125 933.125 -14.795 ;
        RECT 931.435 -15.125 931.765 -14.795 ;
        RECT 930.075 -15.125 930.405 -14.795 ;
        RECT 928.715 -15.125 929.045 -14.795 ;
        RECT 927.355 -15.125 927.685 -14.795 ;
        RECT 925.995 -15.125 926.325 -14.795 ;
        RECT 924.635 -15.125 924.965 -14.795 ;
        RECT 923.275 -15.125 923.605 -14.795 ;
        RECT 921.915 -15.125 922.245 -14.795 ;
        RECT 920.555 -15.125 920.885 -14.795 ;
        RECT 919.195 -15.125 919.525 -14.795 ;
        RECT 917.835 -15.125 918.165 -14.795 ;
        RECT 916.475 -15.125 916.805 -14.795 ;
        RECT 915.115 -15.125 915.445 -14.795 ;
        RECT 913.755 -15.125 914.085 -14.795 ;
        RECT 912.395 -15.125 912.725 -14.795 ;
        RECT 911.035 -15.125 911.365 -14.795 ;
        RECT 909.675 -15.125 910.005 -14.795 ;
        RECT 908.315 -15.125 908.645 -14.795 ;
        RECT 906.955 -15.125 907.285 -14.795 ;
        RECT 905.595 -15.125 905.925 -14.795 ;
        RECT 904.235 -15.125 904.565 -14.795 ;
        RECT 902.875 -15.125 903.205 -14.795 ;
        RECT 901.515 -15.125 901.845 -14.795 ;
        RECT 900.155 -15.125 900.485 -14.795 ;
        RECT 898.795 -15.125 899.125 -14.795 ;
        RECT 897.435 -15.125 897.765 -14.795 ;
        RECT 896.075 -15.125 896.405 -14.795 ;
        RECT 894.715 -15.125 895.045 -14.795 ;
        RECT 893.355 -15.125 893.685 -14.795 ;
        RECT 891.995 -15.125 892.325 -14.795 ;
        RECT 890.635 -15.125 890.965 -14.795 ;
        RECT 889.275 -15.125 889.605 -14.795 ;
        RECT 887.915 -15.125 888.245 -14.795 ;
        RECT 886.555 -15.125 886.885 -14.795 ;
        RECT 885.195 -15.125 885.525 -14.795 ;
        RECT 883.835 -15.125 884.165 -14.795 ;
        RECT 882.475 -15.125 882.805 -14.795 ;
        RECT 881.115 -15.125 881.445 -14.795 ;
        RECT 879.755 -15.125 880.085 -14.795 ;
        RECT 878.395 -15.125 878.725 -14.795 ;
        RECT 877.035 -15.125 877.365 -14.795 ;
        RECT 875.675 -15.125 876.005 -14.795 ;
        RECT 874.315 -15.125 874.645 -14.795 ;
        RECT 872.955 -15.125 873.285 -14.795 ;
        RECT 871.595 -15.125 871.925 -14.795 ;
        RECT 870.235 -15.125 870.565 -14.795 ;
        RECT 868.875 -15.125 869.205 -14.795 ;
        RECT 867.515 -15.125 867.845 -14.795 ;
        RECT 866.155 -15.125 866.485 -14.795 ;
        RECT 864.795 -15.125 865.125 -14.795 ;
        RECT 863.435 -15.125 863.765 -14.795 ;
        RECT 862.075 -15.125 862.405 -14.795 ;
        RECT 860.715 -15.125 861.045 -14.795 ;
        RECT 859.355 -15.125 859.685 -14.795 ;
        RECT 857.995 -15.125 858.325 -14.795 ;
        RECT 856.635 -15.125 856.965 -14.795 ;
        RECT 855.275 -15.125 855.605 -14.795 ;
        RECT 853.915 -15.125 854.245 -14.795 ;
        RECT 852.555 -15.125 852.885 -14.795 ;
        RECT 851.195 -15.125 851.525 -14.795 ;
        RECT 849.835 -15.125 850.165 -14.795 ;
        RECT 848.475 -15.125 848.805 -14.795 ;
        RECT 847.115 -15.125 847.445 -14.795 ;
        RECT 845.755 -15.125 846.085 -14.795 ;
        RECT 844.395 -15.125 844.725 -14.795 ;
        RECT 843.035 -15.125 843.365 -14.795 ;
        RECT 841.675 -15.125 842.005 -14.795 ;
        RECT 840.315 -15.125 840.645 -14.795 ;
        RECT 838.955 -15.125 839.285 -14.795 ;
        RECT 837.595 -15.125 837.925 -14.795 ;
        RECT 836.235 -15.125 836.565 -14.795 ;
        RECT 834.875 -15.125 835.205 -14.795 ;
        RECT 833.515 -15.125 833.845 -14.795 ;
        RECT 832.155 -15.125 832.485 -14.795 ;
        RECT 830.795 -15.125 831.125 -14.795 ;
        RECT 829.435 -15.125 829.765 -14.795 ;
        RECT 828.075 -15.125 828.405 -14.795 ;
        RECT 826.715 -15.125 827.045 -14.795 ;
        RECT 825.355 -15.125 825.685 -14.795 ;
        RECT 823.995 -15.125 824.325 -14.795 ;
        RECT 822.635 -15.125 822.965 -14.795 ;
        RECT 821.275 -15.125 821.605 -14.795 ;
        RECT 819.915 -15.125 820.245 -14.795 ;
        RECT 818.555 -15.125 818.885 -14.795 ;
        RECT 817.195 -15.125 817.525 -14.795 ;
        RECT 815.835 -15.125 816.165 -14.795 ;
        RECT 814.475 -15.125 814.805 -14.795 ;
        RECT 813.115 -15.125 813.445 -14.795 ;
        RECT 811.755 -15.125 812.085 -14.795 ;
        RECT 810.395 -15.125 810.725 -14.795 ;
        RECT 809.035 -15.125 809.365 -14.795 ;
        RECT 807.675 -15.125 808.005 -14.795 ;
        RECT 806.315 -15.125 806.645 -14.795 ;
        RECT 804.955 -15.125 805.285 -14.795 ;
        RECT 803.595 -15.125 803.925 -14.795 ;
        RECT 802.235 -15.125 802.565 -14.795 ;
        RECT 800.875 -15.125 801.205 -14.795 ;
        RECT 799.515 -15.125 799.845 -14.795 ;
        RECT 798.155 -15.125 798.485 -14.795 ;
        RECT 796.795 -15.125 797.125 -14.795 ;
        RECT 795.435 -15.125 795.765 -14.795 ;
        RECT 794.075 -15.125 794.405 -14.795 ;
        RECT 792.715 -15.125 793.045 -14.795 ;
        RECT 791.355 -15.125 791.685 -14.795 ;
        RECT 789.995 -15.125 790.325 -14.795 ;
        RECT 788.635 -15.125 788.965 -14.795 ;
        RECT 787.275 -15.125 787.605 -14.795 ;
        RECT 785.915 -15.125 786.245 -14.795 ;
        RECT 784.555 -15.125 784.885 -14.795 ;
        RECT 783.195 -15.125 783.525 -14.795 ;
        RECT 781.835 -15.125 782.165 -14.795 ;
        RECT 780.475 -15.125 780.805 -14.795 ;
        RECT 779.115 -15.125 779.445 -14.795 ;
        RECT 777.755 -15.125 778.085 -14.795 ;
        RECT 776.395 -15.125 776.725 -14.795 ;
        RECT 775.035 -15.125 775.365 -14.795 ;
        RECT 773.675 -15.125 774.005 -14.795 ;
        RECT 772.315 -15.125 772.645 -14.795 ;
        RECT 770.955 -15.125 771.285 -14.795 ;
        RECT 769.595 -15.125 769.925 -14.795 ;
        RECT 768.235 -15.125 768.565 -14.795 ;
        RECT 766.875 -15.125 767.205 -14.795 ;
        RECT 765.515 -15.125 765.845 -14.795 ;
        RECT 764.155 -15.125 764.485 -14.795 ;
        RECT 762.795 -15.125 763.125 -14.795 ;
        RECT 761.435 -15.125 761.765 -14.795 ;
        RECT 760.075 -15.125 760.405 -14.795 ;
        RECT 758.715 -15.125 759.045 -14.795 ;
        RECT 757.355 -15.125 757.685 -14.795 ;
        RECT 755.995 -15.125 756.325 -14.795 ;
        RECT 754.635 -15.125 754.965 -14.795 ;
        RECT 753.275 -15.125 753.605 -14.795 ;
        RECT 751.915 -15.125 752.245 -14.795 ;
        RECT 750.555 -15.125 750.885 -14.795 ;
        RECT 749.195 -15.125 749.525 -14.795 ;
        RECT 747.835 -15.125 748.165 -14.795 ;
        RECT 746.475 -15.125 746.805 -14.795 ;
        RECT 745.115 -15.125 745.445 -14.795 ;
        RECT 743.755 -15.125 744.085 -14.795 ;
        RECT 742.395 -15.125 742.725 -14.795 ;
        RECT 741.035 -15.125 741.365 -14.795 ;
        RECT 739.675 -15.125 740.005 -14.795 ;
        RECT 738.315 -15.125 738.645 -14.795 ;
        RECT 736.955 -15.125 737.285 -14.795 ;
        RECT 735.595 -15.125 735.925 -14.795 ;
        RECT 734.235 -15.125 734.565 -14.795 ;
        RECT 732.875 -15.125 733.205 -14.795 ;
        RECT 731.515 -15.125 731.845 -14.795 ;
        RECT 730.155 -15.125 730.485 -14.795 ;
        RECT 728.795 -15.125 729.125 -14.795 ;
        RECT 727.435 -15.125 727.765 -14.795 ;
        RECT 726.075 -15.125 726.405 -14.795 ;
        RECT 724.715 -15.125 725.045 -14.795 ;
        RECT 723.355 -15.125 723.685 -14.795 ;
        RECT 721.995 -15.125 722.325 -14.795 ;
        RECT 720.635 -15.125 720.965 -14.795 ;
        RECT 719.275 -15.125 719.605 -14.795 ;
        RECT 717.915 -15.125 718.245 -14.795 ;
        RECT 716.555 -15.125 716.885 -14.795 ;
        RECT 715.195 -15.125 715.525 -14.795 ;
        RECT 713.835 -15.125 714.165 -14.795 ;
        RECT 712.475 -15.125 712.805 -14.795 ;
        RECT 711.115 -15.125 711.445 -14.795 ;
        RECT 709.755 -15.125 710.085 -14.795 ;
        RECT 708.395 -15.125 708.725 -14.795 ;
        RECT 707.035 -15.125 707.365 -14.795 ;
        RECT 705.675 -15.125 706.005 -14.795 ;
        RECT 704.315 -15.125 704.645 -14.795 ;
        RECT 702.955 -15.125 703.285 -14.795 ;
        RECT 701.595 -15.125 701.925 -14.795 ;
        RECT 700.235 -15.125 700.565 -14.795 ;
        RECT 698.875 -15.125 699.205 -14.795 ;
        RECT 697.515 -15.125 697.845 -14.795 ;
        RECT 696.155 -15.125 696.485 -14.795 ;
        RECT 694.795 -15.125 695.125 -14.795 ;
        RECT 693.435 -15.125 693.765 -14.795 ;
        RECT 692.075 -15.125 692.405 -14.795 ;
        RECT 690.715 -15.125 691.045 -14.795 ;
        RECT 689.355 -15.125 689.685 -14.795 ;
        RECT 687.995 -15.125 688.325 -14.795 ;
        RECT 686.635 -15.125 686.965 -14.795 ;
        RECT 685.275 -15.125 685.605 -14.795 ;
        RECT 683.915 -15.125 684.245 -14.795 ;
        RECT 682.555 -15.125 682.885 -14.795 ;
        RECT 681.195 -15.125 681.525 -14.795 ;
        RECT 679.835 -15.125 680.165 -14.795 ;
        RECT 678.475 -15.125 678.805 -14.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.115 -16.485 643.445 -16.155 ;
        RECT 641.755 -16.485 642.085 -16.155 ;
        RECT 640.395 -16.485 640.725 -16.155 ;
        RECT 639.035 -16.485 639.365 -16.155 ;
        RECT 637.675 -16.485 638.005 -16.155 ;
        RECT 636.315 -16.485 636.645 -16.155 ;
        RECT 634.955 -16.485 635.285 -16.155 ;
        RECT 633.595 -16.485 633.925 -16.155 ;
        RECT 632.235 -16.485 632.565 -16.155 ;
        RECT 630.875 -16.485 631.205 -16.155 ;
        RECT 629.515 -16.485 629.845 -16.155 ;
        RECT 628.155 -16.485 628.485 -16.155 ;
        RECT 626.795 -16.485 627.125 -16.155 ;
        RECT 625.435 -16.485 625.765 -16.155 ;
        RECT 624.075 -16.485 624.405 -16.155 ;
        RECT 622.715 -16.485 623.045 -16.155 ;
        RECT 621.355 -16.485 621.685 -16.155 ;
        RECT 619.995 -16.485 620.325 -16.155 ;
        RECT 618.635 -16.485 618.965 -16.155 ;
        RECT 617.275 -16.485 617.605 -16.155 ;
        RECT 615.915 -16.485 616.245 -16.155 ;
        RECT 614.555 -16.485 614.885 -16.155 ;
        RECT 613.195 -16.485 613.525 -16.155 ;
        RECT 611.835 -16.485 612.165 -16.155 ;
        RECT 610.475 -16.485 610.805 -16.155 ;
        RECT 609.115 -16.485 609.445 -16.155 ;
        RECT 607.755 -16.485 608.085 -16.155 ;
        RECT 606.395 -16.485 606.725 -16.155 ;
        RECT 605.035 -16.485 605.365 -16.155 ;
        RECT 603.675 -16.485 604.005 -16.155 ;
        RECT 602.315 -16.485 602.645 -16.155 ;
        RECT 600.955 -16.485 601.285 -16.155 ;
        RECT 599.595 -16.485 599.925 -16.155 ;
        RECT 598.235 -16.485 598.565 -16.155 ;
        RECT 596.875 -16.485 597.205 -16.155 ;
        RECT 595.515 -16.485 595.845 -16.155 ;
        RECT 594.155 -16.485 594.485 -16.155 ;
        RECT 592.795 -16.485 593.125 -16.155 ;
        RECT 591.435 -16.485 591.765 -16.155 ;
        RECT 590.075 -16.485 590.405 -16.155 ;
        RECT 588.715 -16.485 589.045 -16.155 ;
        RECT 587.355 -16.485 587.685 -16.155 ;
        RECT 585.995 -16.485 586.325 -16.155 ;
        RECT 584.635 -16.485 584.965 -16.155 ;
        RECT 583.275 -16.485 583.605 -16.155 ;
        RECT 581.915 -16.485 582.245 -16.155 ;
        RECT 580.555 -16.485 580.885 -16.155 ;
        RECT 579.195 -16.485 579.525 -16.155 ;
        RECT 577.835 -16.485 578.165 -16.155 ;
        RECT 576.475 -16.485 576.805 -16.155 ;
        RECT 575.115 -16.485 575.445 -16.155 ;
        RECT 573.755 -16.485 574.085 -16.155 ;
        RECT 572.395 -16.485 572.725 -16.155 ;
        RECT 571.035 -16.485 571.365 -16.155 ;
        RECT 569.675 -16.485 570.005 -16.155 ;
        RECT 568.315 -16.485 568.645 -16.155 ;
        RECT 566.955 -16.485 567.285 -16.155 ;
        RECT 565.595 -16.485 565.925 -16.155 ;
        RECT 564.235 -16.485 564.565 -16.155 ;
        RECT 562.875 -16.485 563.205 -16.155 ;
        RECT 561.515 -16.485 561.845 -16.155 ;
        RECT 560.155 -16.485 560.485 -16.155 ;
        RECT 558.795 -16.485 559.125 -16.155 ;
        RECT 557.435 -16.485 557.765 -16.155 ;
        RECT 556.075 -16.485 556.405 -16.155 ;
        RECT 554.715 -16.485 555.045 -16.155 ;
        RECT 553.355 -16.485 553.685 -16.155 ;
        RECT 551.995 -16.485 552.325 -16.155 ;
        RECT 550.635 -16.485 550.965 -16.155 ;
        RECT 549.275 -16.485 549.605 -16.155 ;
        RECT 547.915 -16.485 548.245 -16.155 ;
        RECT 546.555 -16.485 546.885 -16.155 ;
        RECT 545.195 -16.485 545.525 -16.155 ;
        RECT 543.835 -16.485 544.165 -16.155 ;
        RECT 542.475 -16.485 542.805 -16.155 ;
        RECT 541.115 -16.485 541.445 -16.155 ;
        RECT 539.755 -16.485 540.085 -16.155 ;
        RECT 538.395 -16.485 538.725 -16.155 ;
        RECT 537.035 -16.485 537.365 -16.155 ;
        RECT 535.675 -16.485 536.005 -16.155 ;
        RECT 534.315 -16.485 534.645 -16.155 ;
        RECT 532.955 -16.485 533.285 -16.155 ;
        RECT 531.595 -16.485 531.925 -16.155 ;
        RECT 530.235 -16.485 530.565 -16.155 ;
        RECT 528.875 -16.485 529.205 -16.155 ;
        RECT 527.515 -16.485 527.845 -16.155 ;
        RECT 526.155 -16.485 526.485 -16.155 ;
        RECT 524.795 -16.485 525.125 -16.155 ;
        RECT 523.435 -16.485 523.765 -16.155 ;
        RECT 522.075 -16.485 522.405 -16.155 ;
        RECT 520.715 -16.485 521.045 -16.155 ;
        RECT 519.355 -16.485 519.685 -16.155 ;
        RECT 517.995 -16.485 518.325 -16.155 ;
        RECT 516.635 -16.485 516.965 -16.155 ;
        RECT 515.275 -16.485 515.605 -16.155 ;
        RECT 513.915 -16.485 514.245 -16.155 ;
        RECT 512.555 -16.485 512.885 -16.155 ;
        RECT 511.195 -16.485 511.525 -16.155 ;
        RECT 509.835 -16.485 510.165 -16.155 ;
        RECT 508.475 -16.485 508.805 -16.155 ;
        RECT 507.115 -16.485 507.445 -16.155 ;
        RECT 505.755 -16.485 506.085 -16.155 ;
        RECT 504.395 -16.485 504.725 -16.155 ;
        RECT 503.035 -16.485 503.365 -16.155 ;
        RECT 501.675 -16.485 502.005 -16.155 ;
        RECT 500.315 -16.485 500.645 -16.155 ;
        RECT 498.955 -16.485 499.285 -16.155 ;
        RECT 497.595 -16.485 497.925 -16.155 ;
        RECT 496.235 -16.485 496.565 -16.155 ;
        RECT 494.875 -16.485 495.205 -16.155 ;
        RECT 493.515 -16.485 493.845 -16.155 ;
        RECT 492.155 -16.485 492.485 -16.155 ;
        RECT 490.795 -16.485 491.125 -16.155 ;
        RECT 489.435 -16.485 489.765 -16.155 ;
        RECT 488.075 -16.485 488.405 -16.155 ;
        RECT 486.715 -16.485 487.045 -16.155 ;
        RECT 485.355 -16.485 485.685 -16.155 ;
        RECT 483.995 -16.485 484.325 -16.155 ;
        RECT 482.635 -16.485 482.965 -16.155 ;
        RECT 481.275 -16.485 481.605 -16.155 ;
        RECT 479.915 -16.485 480.245 -16.155 ;
        RECT 478.555 -16.485 478.885 -16.155 ;
        RECT 477.195 -16.485 477.525 -16.155 ;
        RECT 475.835 -16.485 476.165 -16.155 ;
        RECT 474.475 -16.485 474.805 -16.155 ;
        RECT 473.115 -16.485 473.445 -16.155 ;
        RECT 471.755 -16.485 472.085 -16.155 ;
        RECT 470.395 -16.485 470.725 -16.155 ;
        RECT 469.035 -16.485 469.365 -16.155 ;
        RECT 467.675 -16.485 468.005 -16.155 ;
        RECT 466.315 -16.485 466.645 -16.155 ;
        RECT 464.955 -16.485 465.285 -16.155 ;
        RECT 463.595 -16.485 463.925 -16.155 ;
        RECT 462.235 -16.485 462.565 -16.155 ;
        RECT 460.875 -16.485 461.205 -16.155 ;
        RECT 459.515 -16.485 459.845 -16.155 ;
        RECT 458.155 -16.485 458.485 -16.155 ;
        RECT 456.795 -16.485 457.125 -16.155 ;
        RECT 455.435 -16.485 455.765 -16.155 ;
        RECT 454.075 -16.485 454.405 -16.155 ;
        RECT 452.715 -16.485 453.045 -16.155 ;
        RECT 451.355 -16.485 451.685 -16.155 ;
        RECT 449.995 -16.485 450.325 -16.155 ;
        RECT 448.635 -16.485 448.965 -16.155 ;
        RECT 447.275 -16.485 447.605 -16.155 ;
        RECT 445.915 -16.485 446.245 -16.155 ;
        RECT 444.555 -16.485 444.885 -16.155 ;
        RECT 443.195 -16.485 443.525 -16.155 ;
        RECT 441.835 -16.485 442.165 -16.155 ;
        RECT 440.475 -16.485 440.805 -16.155 ;
        RECT 439.115 -16.485 439.445 -16.155 ;
        RECT 437.755 -16.485 438.085 -16.155 ;
        RECT 436.395 -16.485 436.725 -16.155 ;
        RECT 435.035 -16.485 435.365 -16.155 ;
        RECT 433.675 -16.485 434.005 -16.155 ;
        RECT 432.315 -16.485 432.645 -16.155 ;
        RECT 430.955 -16.485 431.285 -16.155 ;
        RECT 429.595 -16.485 429.925 -16.155 ;
        RECT 428.235 -16.485 428.565 -16.155 ;
        RECT 426.875 -16.485 427.205 -16.155 ;
        RECT 425.515 -16.485 425.845 -16.155 ;
        RECT 424.155 -16.485 424.485 -16.155 ;
        RECT 422.795 -16.485 423.125 -16.155 ;
        RECT 421.435 -16.485 421.765 -16.155 ;
        RECT 420.075 -16.485 420.405 -16.155 ;
        RECT 418.715 -16.485 419.045 -16.155 ;
        RECT 417.355 -16.485 417.685 -16.155 ;
        RECT 415.995 -16.485 416.325 -16.155 ;
        RECT 414.635 -16.485 414.965 -16.155 ;
        RECT 413.275 -16.485 413.605 -16.155 ;
        RECT 411.915 -16.485 412.245 -16.155 ;
        RECT 410.555 -16.485 410.885 -16.155 ;
        RECT 409.195 -16.485 409.525 -16.155 ;
        RECT 407.835 -16.485 408.165 -16.155 ;
        RECT 406.475 -16.485 406.805 -16.155 ;
        RECT 405.115 -16.485 405.445 -16.155 ;
        RECT 403.755 -16.485 404.085 -16.155 ;
        RECT 402.395 -16.485 402.725 -16.155 ;
        RECT 401.035 -16.485 401.365 -16.155 ;
        RECT 399.675 -16.485 400.005 -16.155 ;
        RECT 398.315 -16.485 398.645 -16.155 ;
        RECT 396.955 -16.485 397.285 -16.155 ;
        RECT 395.595 -16.485 395.925 -16.155 ;
        RECT 394.235 -16.485 394.565 -16.155 ;
        RECT 392.875 -16.485 393.205 -16.155 ;
        RECT 391.515 -16.485 391.845 -16.155 ;
        RECT 390.155 -16.485 390.485 -16.155 ;
        RECT 388.795 -16.485 389.125 -16.155 ;
        RECT 387.435 -16.485 387.765 -16.155 ;
        RECT 386.075 -16.485 386.405 -16.155 ;
        RECT 384.715 -16.485 385.045 -16.155 ;
        RECT 383.355 -16.485 383.685 -16.155 ;
        RECT 381.995 -16.485 382.325 -16.155 ;
        RECT 380.635 -16.485 380.965 -16.155 ;
        RECT 379.275 -16.485 379.605 -16.155 ;
        RECT 377.915 -16.485 378.245 -16.155 ;
        RECT 376.555 -16.485 376.885 -16.155 ;
        RECT 375.195 -16.485 375.525 -16.155 ;
        RECT 373.835 -16.485 374.165 -16.155 ;
        RECT 372.475 -16.485 372.805 -16.155 ;
        RECT 371.115 -16.485 371.445 -16.155 ;
        RECT 369.755 -16.485 370.085 -16.155 ;
        RECT 368.395 -16.485 368.725 -16.155 ;
        RECT 367.035 -16.485 367.365 -16.155 ;
        RECT 365.675 -16.485 366.005 -16.155 ;
        RECT 364.315 -16.485 364.645 -16.155 ;
        RECT 362.955 -16.485 363.285 -16.155 ;
        RECT 361.595 -16.485 361.925 -16.155 ;
        RECT 360.235 -16.485 360.565 -16.155 ;
        RECT 358.875 -16.485 359.205 -16.155 ;
        RECT 357.515 -16.485 357.845 -16.155 ;
        RECT 356.155 -16.485 356.485 -16.155 ;
        RECT 354.795 -16.485 355.125 -16.155 ;
        RECT 353.435 -16.485 353.765 -16.155 ;
        RECT 352.075 -16.485 352.405 -16.155 ;
        RECT 350.715 -16.485 351.045 -16.155 ;
        RECT 349.355 -16.485 349.685 -16.155 ;
        RECT 347.995 -16.485 348.325 -16.155 ;
        RECT 346.635 -16.485 346.965 -16.155 ;
        RECT 345.275 -16.485 345.605 -16.155 ;
        RECT 343.915 -16.485 344.245 -16.155 ;
        RECT 342.555 -16.485 342.885 -16.155 ;
        RECT 341.195 -16.485 341.525 -16.155 ;
        RECT 339.835 -16.485 340.165 -16.155 ;
        RECT 338.475 -16.485 338.805 -16.155 ;
        RECT 337.115 -16.485 337.445 -16.155 ;
        RECT 335.755 -16.485 336.085 -16.155 ;
        RECT 334.395 -16.485 334.725 -16.155 ;
        RECT 333.035 -16.485 333.365 -16.155 ;
        RECT 331.675 -16.485 332.005 -16.155 ;
        RECT 330.315 -16.485 330.645 -16.155 ;
        RECT 328.955 -16.485 329.285 -16.155 ;
        RECT 327.595 -16.485 327.925 -16.155 ;
        RECT 326.235 -16.485 326.565 -16.155 ;
        RECT 324.875 -16.485 325.205 -16.155 ;
        RECT 323.515 -16.485 323.845 -16.155 ;
        RECT 322.155 -16.485 322.485 -16.155 ;
        RECT 320.795 -16.485 321.125 -16.155 ;
        RECT 319.435 -16.485 319.765 -16.155 ;
        RECT 318.075 -16.485 318.405 -16.155 ;
        RECT 316.715 -16.485 317.045 -16.155 ;
        RECT 315.355 -16.485 315.685 -16.155 ;
        RECT 313.995 -16.485 314.325 -16.155 ;
        RECT 312.635 -16.485 312.965 -16.155 ;
        RECT 311.275 -16.485 311.605 -16.155 ;
        RECT 309.915 -16.485 310.245 -16.155 ;
        RECT 308.555 -16.485 308.885 -16.155 ;
        RECT 307.195 -16.485 307.525 -16.155 ;
        RECT 305.835 -16.485 306.165 -16.155 ;
        RECT 304.475 -16.485 304.805 -16.155 ;
        RECT 303.115 -16.485 303.445 -16.155 ;
        RECT 301.755 -16.485 302.085 -16.155 ;
        RECT 300.395 -16.485 300.725 -16.155 ;
        RECT 299.035 -16.485 299.365 -16.155 ;
        RECT 297.675 -16.485 298.005 -16.155 ;
        RECT 296.315 -16.485 296.645 -16.155 ;
        RECT 294.955 -16.485 295.285 -16.155 ;
        RECT 293.595 -16.485 293.925 -16.155 ;
        RECT 292.235 -16.485 292.565 -16.155 ;
        RECT 290.875 -16.485 291.205 -16.155 ;
        RECT 289.515 -16.485 289.845 -16.155 ;
        RECT 288.155 -16.485 288.485 -16.155 ;
        RECT 286.795 -16.485 287.125 -16.155 ;
        RECT 285.435 -16.485 285.765 -16.155 ;
        RECT 284.075 -16.485 284.405 -16.155 ;
        RECT 282.715 -16.485 283.045 -16.155 ;
        RECT 281.355 -16.485 281.685 -16.155 ;
        RECT 279.995 -16.485 280.325 -16.155 ;
        RECT 278.635 -16.485 278.965 -16.155 ;
        RECT 277.275 -16.485 277.605 -16.155 ;
        RECT 275.915 -16.485 276.245 -16.155 ;
        RECT 274.555 -16.485 274.885 -16.155 ;
        RECT 273.195 -16.485 273.525 -16.155 ;
        RECT 271.835 -16.485 272.165 -16.155 ;
        RECT 270.475 -16.485 270.805 -16.155 ;
        RECT 269.115 -16.485 269.445 -16.155 ;
        RECT 267.755 -16.485 268.085 -16.155 ;
        RECT 266.395 -16.485 266.725 -16.155 ;
        RECT 265.035 -16.485 265.365 -16.155 ;
        RECT 263.675 -16.485 264.005 -16.155 ;
        RECT 262.315 -16.485 262.645 -16.155 ;
        RECT 260.955 -16.485 261.285 -16.155 ;
        RECT 259.595 -16.485 259.925 -16.155 ;
        RECT 258.235 -16.485 258.565 -16.155 ;
        RECT 256.875 -16.485 257.205 -16.155 ;
        RECT 255.515 -16.485 255.845 -16.155 ;
        RECT 254.155 -16.485 254.485 -16.155 ;
        RECT 252.795 -16.485 253.125 -16.155 ;
        RECT 251.435 -16.485 251.765 -16.155 ;
        RECT 250.075 -16.485 250.405 -16.155 ;
        RECT 248.715 -16.485 249.045 -16.155 ;
        RECT 247.355 -16.485 247.685 -16.155 ;
        RECT 245.995 -16.485 246.325 -16.155 ;
        RECT 244.635 -16.485 244.965 -16.155 ;
        RECT 243.275 -16.485 243.605 -16.155 ;
        RECT 241.915 -16.485 242.245 -16.155 ;
        RECT 240.555 -16.485 240.885 -16.155 ;
        RECT 239.195 -16.485 239.525 -16.155 ;
        RECT 237.835 -16.485 238.165 -16.155 ;
        RECT 236.475 -16.485 236.805 -16.155 ;
        RECT 235.115 -16.485 235.445 -16.155 ;
        RECT 233.755 -16.485 234.085 -16.155 ;
        RECT 232.395 -16.485 232.725 -16.155 ;
        RECT 231.035 -16.485 231.365 -16.155 ;
        RECT 229.675 -16.485 230.005 -16.155 ;
        RECT 228.315 -16.485 228.645 -16.155 ;
        RECT 226.955 -16.485 227.285 -16.155 ;
        RECT 225.595 -16.485 225.925 -16.155 ;
        RECT 224.235 -16.485 224.565 -16.155 ;
        RECT 222.875 -16.485 223.205 -16.155 ;
        RECT 221.515 -16.485 221.845 -16.155 ;
        RECT 220.155 -16.485 220.485 -16.155 ;
        RECT 218.795 -16.485 219.125 -16.155 ;
        RECT 217.435 -16.485 217.765 -16.155 ;
        RECT 216.075 -16.485 216.405 -16.155 ;
        RECT 214.715 -16.485 215.045 -16.155 ;
        RECT 213.355 -16.485 213.685 -16.155 ;
        RECT 211.995 -16.485 212.325 -16.155 ;
        RECT 210.635 -16.485 210.965 -16.155 ;
        RECT 209.275 -16.485 209.605 -16.155 ;
        RECT 207.915 -16.485 208.245 -16.155 ;
        RECT 206.555 -16.485 206.885 -16.155 ;
        RECT 205.195 -16.485 205.525 -16.155 ;
        RECT 203.835 -16.485 204.165 -16.155 ;
        RECT 202.475 -16.485 202.805 -16.155 ;
        RECT 201.115 -16.485 201.445 -16.155 ;
        RECT 199.755 -16.485 200.085 -16.155 ;
        RECT 198.395 -16.485 198.725 -16.155 ;
        RECT 197.035 -16.485 197.365 -16.155 ;
        RECT 195.675 -16.485 196.005 -16.155 ;
        RECT 194.315 -16.485 194.645 -16.155 ;
        RECT 192.955 -16.485 193.285 -16.155 ;
        RECT 191.595 -16.485 191.925 -16.155 ;
        RECT 190.235 -16.485 190.565 -16.155 ;
        RECT 188.875 -16.485 189.205 -16.155 ;
        RECT 187.515 -16.485 187.845 -16.155 ;
        RECT 186.155 -16.485 186.485 -16.155 ;
        RECT 184.795 -16.485 185.125 -16.155 ;
        RECT 183.435 -16.485 183.765 -16.155 ;
        RECT 182.075 -16.485 182.405 -16.155 ;
        RECT 180.715 -16.485 181.045 -16.155 ;
        RECT 179.355 -16.485 179.685 -16.155 ;
        RECT 177.995 -16.485 178.325 -16.155 ;
        RECT 176.635 -16.485 176.965 -16.155 ;
        RECT 175.275 -16.485 175.605 -16.155 ;
        RECT 173.915 -16.485 174.245 -16.155 ;
        RECT 172.555 -16.485 172.885 -16.155 ;
        RECT 171.195 -16.485 171.525 -16.155 ;
        RECT 169.835 -16.485 170.165 -16.155 ;
        RECT 168.475 -16.485 168.805 -16.155 ;
        RECT 167.115 -16.485 167.445 -16.155 ;
        RECT 165.755 -16.485 166.085 -16.155 ;
        RECT 164.395 -16.485 164.725 -16.155 ;
        RECT 163.035 -16.485 163.365 -16.155 ;
        RECT 161.675 -16.485 162.005 -16.155 ;
        RECT 160.315 -16.485 160.645 -16.155 ;
        RECT 158.955 -16.485 159.285 -16.155 ;
        RECT 157.595 -16.485 157.925 -16.155 ;
        RECT 156.235 -16.485 156.565 -16.155 ;
        RECT 154.875 -16.485 155.205 -16.155 ;
        RECT 153.515 -16.485 153.845 -16.155 ;
        RECT 152.155 -16.485 152.485 -16.155 ;
        RECT 150.795 -16.485 151.125 -16.155 ;
        RECT 149.435 -16.485 149.765 -16.155 ;
        RECT 148.075 -16.485 148.405 -16.155 ;
        RECT 146.715 -16.485 147.045 -16.155 ;
        RECT 145.355 -16.485 145.685 -16.155 ;
        RECT 143.995 -16.485 144.325 -16.155 ;
        RECT 142.635 -16.485 142.965 -16.155 ;
        RECT 141.275 -16.485 141.605 -16.155 ;
        RECT 139.915 -16.485 140.245 -16.155 ;
        RECT 138.555 -16.485 138.885 -16.155 ;
        RECT 137.195 -16.485 137.525 -16.155 ;
        RECT 135.835 -16.485 136.165 -16.155 ;
        RECT 134.475 -16.485 134.805 -16.155 ;
        RECT 133.115 -16.485 133.445 -16.155 ;
        RECT 131.755 -16.485 132.085 -16.155 ;
        RECT 130.395 -16.485 130.725 -16.155 ;
        RECT 129.035 -16.485 129.365 -16.155 ;
        RECT 127.675 -16.485 128.005 -16.155 ;
        RECT 126.315 -16.485 126.645 -16.155 ;
        RECT 124.955 -16.485 125.285 -16.155 ;
        RECT 123.595 -16.485 123.925 -16.155 ;
        RECT 122.235 -16.485 122.565 -16.155 ;
        RECT 120.875 -16.485 121.205 -16.155 ;
        RECT 119.515 -16.485 119.845 -16.155 ;
        RECT 118.155 -16.485 118.485 -16.155 ;
        RECT 116.795 -16.485 117.125 -16.155 ;
        RECT 115.435 -16.485 115.765 -16.155 ;
        RECT 114.075 -16.485 114.405 -16.155 ;
        RECT 112.715 -16.485 113.045 -16.155 ;
        RECT 111.355 -16.485 111.685 -16.155 ;
        RECT 109.995 -16.485 110.325 -16.155 ;
        RECT 108.635 -16.485 108.965 -16.155 ;
        RECT 107.275 -16.485 107.605 -16.155 ;
        RECT 105.915 -16.485 106.245 -16.155 ;
        RECT 104.555 -16.485 104.885 -16.155 ;
        RECT 103.195 -16.485 103.525 -16.155 ;
        RECT 101.835 -16.485 102.165 -16.155 ;
        RECT 100.475 -16.485 100.805 -16.155 ;
        RECT 99.115 -16.485 99.445 -16.155 ;
        RECT 97.755 -16.485 98.085 -16.155 ;
        RECT 96.395 -16.485 96.725 -16.155 ;
        RECT 95.035 -16.485 95.365 -16.155 ;
        RECT 93.675 -16.485 94.005 -16.155 ;
        RECT 92.315 -16.485 92.645 -16.155 ;
        RECT 90.955 -16.485 91.285 -16.155 ;
        RECT 89.595 -16.485 89.925 -16.155 ;
        RECT 88.235 -16.485 88.565 -16.155 ;
        RECT 86.875 -16.485 87.205 -16.155 ;
        RECT 85.515 -16.485 85.845 -16.155 ;
        RECT 84.155 -16.485 84.485 -16.155 ;
        RECT 82.795 -16.485 83.125 -16.155 ;
        RECT 81.435 -16.485 81.765 -16.155 ;
        RECT 80.075 -16.485 80.405 -16.155 ;
        RECT 78.715 -16.485 79.045 -16.155 ;
        RECT 77.355 -16.485 77.685 -16.155 ;
        RECT 75.995 -16.485 76.325 -16.155 ;
        RECT 74.635 -16.485 74.965 -16.155 ;
        RECT 73.275 -16.485 73.605 -16.155 ;
        RECT 71.915 -16.485 72.245 -16.155 ;
        RECT 70.555 -16.485 70.885 -16.155 ;
        RECT 69.195 -16.485 69.525 -16.155 ;
        RECT 67.835 -16.485 68.165 -16.155 ;
        RECT 66.475 -16.485 66.805 -16.155 ;
        RECT 65.115 -16.485 65.445 -16.155 ;
        RECT 63.755 -16.485 64.085 -16.155 ;
        RECT 62.395 -16.485 62.725 -16.155 ;
        RECT 61.035 -16.485 61.365 -16.155 ;
        RECT 59.675 -16.485 60.005 -16.155 ;
        RECT 58.315 -16.485 58.645 -16.155 ;
        RECT 56.955 -16.485 57.285 -16.155 ;
        RECT 55.595 -16.485 55.925 -16.155 ;
        RECT 54.235 -16.485 54.565 -16.155 ;
        RECT 52.875 -16.485 53.205 -16.155 ;
        RECT 51.515 -16.485 51.845 -16.155 ;
        RECT 50.155 -16.485 50.485 -16.155 ;
        RECT 48.795 -16.485 49.125 -16.155 ;
        RECT 47.435 -16.485 47.765 -16.155 ;
        RECT 46.075 -16.485 46.405 -16.155 ;
        RECT 44.715 -16.485 45.045 -16.155 ;
        RECT 43.355 -16.485 43.685 -16.155 ;
        RECT 41.995 -16.485 42.325 -16.155 ;
        RECT 40.635 -16.485 40.965 -16.155 ;
        RECT 39.275 -16.485 39.605 -16.155 ;
        RECT 37.915 -16.485 38.245 -16.155 ;
        RECT 36.555 -16.485 36.885 -16.155 ;
        RECT 35.195 -16.485 35.525 -16.155 ;
        RECT 33.835 -16.485 34.165 -16.155 ;
        RECT 32.475 -16.485 32.805 -16.155 ;
        RECT 31.115 -16.485 31.445 -16.155 ;
        RECT 29.755 -16.485 30.085 -16.155 ;
        RECT 28.395 -16.485 28.725 -16.155 ;
        RECT 27.035 -16.485 27.365 -16.155 ;
        RECT 25.675 -16.485 26.005 -16.155 ;
        RECT 24.315 -16.485 24.645 -16.155 ;
        RECT 22.955 -16.485 23.285 -16.155 ;
        RECT 21.595 -16.485 21.925 -16.155 ;
        RECT 20.235 -16.485 20.565 -16.155 ;
        RECT 18.875 -16.485 19.205 -16.155 ;
        RECT 17.515 -16.485 17.845 -16.155 ;
        RECT 16.155 -16.485 16.485 -16.155 ;
        RECT 14.795 -16.485 15.125 -16.155 ;
        RECT 13.435 -16.485 13.765 -16.155 ;
        RECT 12.075 -16.485 12.405 -16.155 ;
        RECT 10.715 -16.485 11.045 -16.155 ;
        RECT 9.355 -16.485 9.685 -16.155 ;
        RECT 7.995 -16.485 8.325 -16.155 ;
        RECT 6.635 -16.485 6.965 -16.155 ;
        RECT 5.275 -16.485 5.605 -16.155 ;
        RECT 3.915 -16.485 4.245 -16.155 ;
        RECT 2.555 -16.485 2.885 -16.155 ;
        RECT 1.195 -16.485 1.525 -16.155 ;
        RECT -0.165 -16.485 0.165 -16.155 ;
        RECT -1.525 -16.485 -1.195 -16.155 ;
        RECT -1.525 -16.48 678.475 -16.16 ;
        RECT 677.115 -16.485 677.445 -16.155 ;
        RECT 675.755 -16.485 676.085 -16.155 ;
        RECT 674.395 -16.485 674.725 -16.155 ;
        RECT 673.035 -16.485 673.365 -16.155 ;
        RECT 671.675 -16.485 672.005 -16.155 ;
        RECT 670.315 -16.485 670.645 -16.155 ;
        RECT 668.955 -16.485 669.285 -16.155 ;
        RECT 667.595 -16.485 667.925 -16.155 ;
        RECT 666.235 -16.485 666.565 -16.155 ;
        RECT 664.875 -16.485 665.205 -16.155 ;
        RECT 663.515 -16.485 663.845 -16.155 ;
        RECT 662.155 -16.485 662.485 -16.155 ;
        RECT 660.795 -16.485 661.125 -16.155 ;
        RECT 659.435 -16.485 659.765 -16.155 ;
        RECT 658.075 -16.485 658.405 -16.155 ;
        RECT 656.715 -16.485 657.045 -16.155 ;
        RECT 655.355 -16.485 655.685 -16.155 ;
        RECT 653.995 -16.485 654.325 -16.155 ;
        RECT 652.635 -16.485 652.965 -16.155 ;
        RECT 651.275 -16.485 651.605 -16.155 ;
        RECT 649.915 -16.485 650.245 -16.155 ;
        RECT 648.555 -16.485 648.885 -16.155 ;
        RECT 647.195 -16.485 647.525 -16.155 ;
        RECT 645.835 -16.485 646.165 -16.155 ;
        RECT 644.475 -16.485 644.805 -16.155 ;
        RECT 954.555 -16.485 954.885 -16.155 ;
        RECT 678.475 -16.48 954.885 -16.16 ;
        RECT 953.195 -16.485 953.525 -16.155 ;
        RECT 951.835 -16.485 952.165 -16.155 ;
        RECT 950.475 -16.485 950.805 -16.155 ;
        RECT 949.115 -16.485 949.445 -16.155 ;
        RECT 947.755 -16.485 948.085 -16.155 ;
        RECT 946.395 -16.485 946.725 -16.155 ;
        RECT 945.035 -16.485 945.365 -16.155 ;
        RECT 943.675 -16.485 944.005 -16.155 ;
        RECT 942.315 -16.485 942.645 -16.155 ;
        RECT 940.955 -16.485 941.285 -16.155 ;
        RECT 939.595 -16.485 939.925 -16.155 ;
        RECT 938.235 -16.485 938.565 -16.155 ;
        RECT 936.875 -16.485 937.205 -16.155 ;
        RECT 935.515 -16.485 935.845 -16.155 ;
        RECT 934.155 -16.485 934.485 -16.155 ;
        RECT 932.795 -16.485 933.125 -16.155 ;
        RECT 931.435 -16.485 931.765 -16.155 ;
        RECT 930.075 -16.485 930.405 -16.155 ;
        RECT 928.715 -16.485 929.045 -16.155 ;
        RECT 927.355 -16.485 927.685 -16.155 ;
        RECT 925.995 -16.485 926.325 -16.155 ;
        RECT 924.635 -16.485 924.965 -16.155 ;
        RECT 923.275 -16.485 923.605 -16.155 ;
        RECT 921.915 -16.485 922.245 -16.155 ;
        RECT 920.555 -16.485 920.885 -16.155 ;
        RECT 919.195 -16.485 919.525 -16.155 ;
        RECT 917.835 -16.485 918.165 -16.155 ;
        RECT 916.475 -16.485 916.805 -16.155 ;
        RECT 915.115 -16.485 915.445 -16.155 ;
        RECT 913.755 -16.485 914.085 -16.155 ;
        RECT 912.395 -16.485 912.725 -16.155 ;
        RECT 911.035 -16.485 911.365 -16.155 ;
        RECT 909.675 -16.485 910.005 -16.155 ;
        RECT 908.315 -16.485 908.645 -16.155 ;
        RECT 906.955 -16.485 907.285 -16.155 ;
        RECT 905.595 -16.485 905.925 -16.155 ;
        RECT 904.235 -16.485 904.565 -16.155 ;
        RECT 902.875 -16.485 903.205 -16.155 ;
        RECT 901.515 -16.485 901.845 -16.155 ;
        RECT 900.155 -16.485 900.485 -16.155 ;
        RECT 898.795 -16.485 899.125 -16.155 ;
        RECT 897.435 -16.485 897.765 -16.155 ;
        RECT 896.075 -16.485 896.405 -16.155 ;
        RECT 894.715 -16.485 895.045 -16.155 ;
        RECT 893.355 -16.485 893.685 -16.155 ;
        RECT 891.995 -16.485 892.325 -16.155 ;
        RECT 890.635 -16.485 890.965 -16.155 ;
        RECT 889.275 -16.485 889.605 -16.155 ;
        RECT 887.915 -16.485 888.245 -16.155 ;
        RECT 886.555 -16.485 886.885 -16.155 ;
        RECT 885.195 -16.485 885.525 -16.155 ;
        RECT 883.835 -16.485 884.165 -16.155 ;
        RECT 882.475 -16.485 882.805 -16.155 ;
        RECT 881.115 -16.485 881.445 -16.155 ;
        RECT 879.755 -16.485 880.085 -16.155 ;
        RECT 878.395 -16.485 878.725 -16.155 ;
        RECT 877.035 -16.485 877.365 -16.155 ;
        RECT 875.675 -16.485 876.005 -16.155 ;
        RECT 874.315 -16.485 874.645 -16.155 ;
        RECT 872.955 -16.485 873.285 -16.155 ;
        RECT 871.595 -16.485 871.925 -16.155 ;
        RECT 870.235 -16.485 870.565 -16.155 ;
        RECT 868.875 -16.485 869.205 -16.155 ;
        RECT 867.515 -16.485 867.845 -16.155 ;
        RECT 866.155 -16.485 866.485 -16.155 ;
        RECT 864.795 -16.485 865.125 -16.155 ;
        RECT 863.435 -16.485 863.765 -16.155 ;
        RECT 862.075 -16.485 862.405 -16.155 ;
        RECT 860.715 -16.485 861.045 -16.155 ;
        RECT 859.355 -16.485 859.685 -16.155 ;
        RECT 857.995 -16.485 858.325 -16.155 ;
        RECT 856.635 -16.485 856.965 -16.155 ;
        RECT 855.275 -16.485 855.605 -16.155 ;
        RECT 853.915 -16.485 854.245 -16.155 ;
        RECT 852.555 -16.485 852.885 -16.155 ;
        RECT 851.195 -16.485 851.525 -16.155 ;
        RECT 849.835 -16.485 850.165 -16.155 ;
        RECT 848.475 -16.485 848.805 -16.155 ;
        RECT 847.115 -16.485 847.445 -16.155 ;
        RECT 845.755 -16.485 846.085 -16.155 ;
        RECT 844.395 -16.485 844.725 -16.155 ;
        RECT 843.035 -16.485 843.365 -16.155 ;
        RECT 841.675 -16.485 842.005 -16.155 ;
        RECT 840.315 -16.485 840.645 -16.155 ;
        RECT 838.955 -16.485 839.285 -16.155 ;
        RECT 837.595 -16.485 837.925 -16.155 ;
        RECT 836.235 -16.485 836.565 -16.155 ;
        RECT 834.875 -16.485 835.205 -16.155 ;
        RECT 833.515 -16.485 833.845 -16.155 ;
        RECT 832.155 -16.485 832.485 -16.155 ;
        RECT 830.795 -16.485 831.125 -16.155 ;
        RECT 829.435 -16.485 829.765 -16.155 ;
        RECT 828.075 -16.485 828.405 -16.155 ;
        RECT 826.715 -16.485 827.045 -16.155 ;
        RECT 825.355 -16.485 825.685 -16.155 ;
        RECT 823.995 -16.485 824.325 -16.155 ;
        RECT 822.635 -16.485 822.965 -16.155 ;
        RECT 821.275 -16.485 821.605 -16.155 ;
        RECT 819.915 -16.485 820.245 -16.155 ;
        RECT 818.555 -16.485 818.885 -16.155 ;
        RECT 817.195 -16.485 817.525 -16.155 ;
        RECT 815.835 -16.485 816.165 -16.155 ;
        RECT 814.475 -16.485 814.805 -16.155 ;
        RECT 813.115 -16.485 813.445 -16.155 ;
        RECT 811.755 -16.485 812.085 -16.155 ;
        RECT 810.395 -16.485 810.725 -16.155 ;
        RECT 809.035 -16.485 809.365 -16.155 ;
        RECT 807.675 -16.485 808.005 -16.155 ;
        RECT 806.315 -16.485 806.645 -16.155 ;
        RECT 804.955 -16.485 805.285 -16.155 ;
        RECT 803.595 -16.485 803.925 -16.155 ;
        RECT 802.235 -16.485 802.565 -16.155 ;
        RECT 800.875 -16.485 801.205 -16.155 ;
        RECT 799.515 -16.485 799.845 -16.155 ;
        RECT 798.155 -16.485 798.485 -16.155 ;
        RECT 796.795 -16.485 797.125 -16.155 ;
        RECT 795.435 -16.485 795.765 -16.155 ;
        RECT 794.075 -16.485 794.405 -16.155 ;
        RECT 792.715 -16.485 793.045 -16.155 ;
        RECT 791.355 -16.485 791.685 -16.155 ;
        RECT 789.995 -16.485 790.325 -16.155 ;
        RECT 788.635 -16.485 788.965 -16.155 ;
        RECT 787.275 -16.485 787.605 -16.155 ;
        RECT 785.915 -16.485 786.245 -16.155 ;
        RECT 784.555 -16.485 784.885 -16.155 ;
        RECT 783.195 -16.485 783.525 -16.155 ;
        RECT 781.835 -16.485 782.165 -16.155 ;
        RECT 780.475 -16.485 780.805 -16.155 ;
        RECT 779.115 -16.485 779.445 -16.155 ;
        RECT 777.755 -16.485 778.085 -16.155 ;
        RECT 776.395 -16.485 776.725 -16.155 ;
        RECT 775.035 -16.485 775.365 -16.155 ;
        RECT 773.675 -16.485 774.005 -16.155 ;
        RECT 772.315 -16.485 772.645 -16.155 ;
        RECT 770.955 -16.485 771.285 -16.155 ;
        RECT 769.595 -16.485 769.925 -16.155 ;
        RECT 768.235 -16.485 768.565 -16.155 ;
        RECT 766.875 -16.485 767.205 -16.155 ;
        RECT 765.515 -16.485 765.845 -16.155 ;
        RECT 764.155 -16.485 764.485 -16.155 ;
        RECT 762.795 -16.485 763.125 -16.155 ;
        RECT 761.435 -16.485 761.765 -16.155 ;
        RECT 760.075 -16.485 760.405 -16.155 ;
        RECT 758.715 -16.485 759.045 -16.155 ;
        RECT 757.355 -16.485 757.685 -16.155 ;
        RECT 755.995 -16.485 756.325 -16.155 ;
        RECT 754.635 -16.485 754.965 -16.155 ;
        RECT 753.275 -16.485 753.605 -16.155 ;
        RECT 751.915 -16.485 752.245 -16.155 ;
        RECT 750.555 -16.485 750.885 -16.155 ;
        RECT 749.195 -16.485 749.525 -16.155 ;
        RECT 747.835 -16.485 748.165 -16.155 ;
        RECT 746.475 -16.485 746.805 -16.155 ;
        RECT 745.115 -16.485 745.445 -16.155 ;
        RECT 743.755 -16.485 744.085 -16.155 ;
        RECT 742.395 -16.485 742.725 -16.155 ;
        RECT 741.035 -16.485 741.365 -16.155 ;
        RECT 739.675 -16.485 740.005 -16.155 ;
        RECT 738.315 -16.485 738.645 -16.155 ;
        RECT 736.955 -16.485 737.285 -16.155 ;
        RECT 735.595 -16.485 735.925 -16.155 ;
        RECT 734.235 -16.485 734.565 -16.155 ;
        RECT 732.875 -16.485 733.205 -16.155 ;
        RECT 731.515 -16.485 731.845 -16.155 ;
        RECT 730.155 -16.485 730.485 -16.155 ;
        RECT 728.795 -16.485 729.125 -16.155 ;
        RECT 727.435 -16.485 727.765 -16.155 ;
        RECT 726.075 -16.485 726.405 -16.155 ;
        RECT 724.715 -16.485 725.045 -16.155 ;
        RECT 723.355 -16.485 723.685 -16.155 ;
        RECT 721.995 -16.485 722.325 -16.155 ;
        RECT 720.635 -16.485 720.965 -16.155 ;
        RECT 719.275 -16.485 719.605 -16.155 ;
        RECT 717.915 -16.485 718.245 -16.155 ;
        RECT 716.555 -16.485 716.885 -16.155 ;
        RECT 715.195 -16.485 715.525 -16.155 ;
        RECT 713.835 -16.485 714.165 -16.155 ;
        RECT 712.475 -16.485 712.805 -16.155 ;
        RECT 711.115 -16.485 711.445 -16.155 ;
        RECT 709.755 -16.485 710.085 -16.155 ;
        RECT 708.395 -16.485 708.725 -16.155 ;
        RECT 707.035 -16.485 707.365 -16.155 ;
        RECT 705.675 -16.485 706.005 -16.155 ;
        RECT 704.315 -16.485 704.645 -16.155 ;
        RECT 702.955 -16.485 703.285 -16.155 ;
        RECT 701.595 -16.485 701.925 -16.155 ;
        RECT 700.235 -16.485 700.565 -16.155 ;
        RECT 698.875 -16.485 699.205 -16.155 ;
        RECT 697.515 -16.485 697.845 -16.155 ;
        RECT 696.155 -16.485 696.485 -16.155 ;
        RECT 694.795 -16.485 695.125 -16.155 ;
        RECT 693.435 -16.485 693.765 -16.155 ;
        RECT 692.075 -16.485 692.405 -16.155 ;
        RECT 690.715 -16.485 691.045 -16.155 ;
        RECT 689.355 -16.485 689.685 -16.155 ;
        RECT 687.995 -16.485 688.325 -16.155 ;
        RECT 686.635 -16.485 686.965 -16.155 ;
        RECT 685.275 -16.485 685.605 -16.155 ;
        RECT 683.915 -16.485 684.245 -16.155 ;
        RECT 682.555 -16.485 682.885 -16.155 ;
        RECT 681.195 -16.485 681.525 -16.155 ;
        RECT 679.835 -16.485 680.165 -16.155 ;
        RECT 678.475 -16.485 678.805 -16.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -12.4 678.475 -12.08 ;
        RECT 677.115 -12.405 677.445 -12.075 ;
        RECT 675.755 -12.405 676.085 -12.075 ;
        RECT 674.395 -12.405 674.725 -12.075 ;
        RECT 673.035 -12.405 673.365 -12.075 ;
        RECT 671.675 -12.405 672.005 -12.075 ;
        RECT 670.315 -12.405 670.645 -12.075 ;
        RECT 668.955 -12.405 669.285 -12.075 ;
        RECT 667.595 -12.405 667.925 -12.075 ;
        RECT 666.235 -12.405 666.565 -12.075 ;
        RECT 664.875 -12.405 665.205 -12.075 ;
        RECT 663.515 -12.405 663.845 -12.075 ;
        RECT 662.155 -12.405 662.485 -12.075 ;
        RECT 660.795 -12.405 661.125 -12.075 ;
        RECT 659.435 -12.405 659.765 -12.075 ;
        RECT 658.075 -12.405 658.405 -12.075 ;
        RECT 656.715 -12.405 657.045 -12.075 ;
        RECT 655.355 -12.405 655.685 -12.075 ;
        RECT 653.995 -12.405 654.325 -12.075 ;
        RECT 652.635 -12.405 652.965 -12.075 ;
        RECT 651.275 -12.405 651.605 -12.075 ;
        RECT 649.915 -12.405 650.245 -12.075 ;
        RECT 648.555 -12.405 648.885 -12.075 ;
        RECT 647.195 -12.405 647.525 -12.075 ;
        RECT 645.835 -12.405 646.165 -12.075 ;
        RECT 644.475 -12.405 644.805 -12.075 ;
        RECT 643.115 -12.405 643.445 -12.075 ;
        RECT 641.755 -12.405 642.085 -12.075 ;
        RECT 640.395 -12.405 640.725 -12.075 ;
        RECT 639.035 -12.405 639.365 -12.075 ;
        RECT 637.675 -12.405 638.005 -12.075 ;
        RECT 636.315 -12.405 636.645 -12.075 ;
        RECT 634.955 -12.405 635.285 -12.075 ;
        RECT 633.595 -12.405 633.925 -12.075 ;
        RECT 632.235 -12.405 632.565 -12.075 ;
        RECT 630.875 -12.405 631.205 -12.075 ;
        RECT 629.515 -12.405 629.845 -12.075 ;
        RECT 628.155 -12.405 628.485 -12.075 ;
        RECT 626.795 -12.405 627.125 -12.075 ;
        RECT 625.435 -12.405 625.765 -12.075 ;
        RECT 624.075 -12.405 624.405 -12.075 ;
        RECT 622.715 -12.405 623.045 -12.075 ;
        RECT 621.355 -12.405 621.685 -12.075 ;
        RECT 619.995 -12.405 620.325 -12.075 ;
        RECT 618.635 -12.405 618.965 -12.075 ;
        RECT 617.275 -12.405 617.605 -12.075 ;
        RECT 615.915 -12.405 616.245 -12.075 ;
        RECT 614.555 -12.405 614.885 -12.075 ;
        RECT 613.195 -12.405 613.525 -12.075 ;
        RECT 611.835 -12.405 612.165 -12.075 ;
        RECT 610.475 -12.405 610.805 -12.075 ;
        RECT 609.115 -12.405 609.445 -12.075 ;
        RECT 607.755 -12.405 608.085 -12.075 ;
        RECT 606.395 -12.405 606.725 -12.075 ;
        RECT 605.035 -12.405 605.365 -12.075 ;
        RECT 603.675 -12.405 604.005 -12.075 ;
        RECT 602.315 -12.405 602.645 -12.075 ;
        RECT 600.955 -12.405 601.285 -12.075 ;
        RECT 599.595 -12.405 599.925 -12.075 ;
        RECT 598.235 -12.405 598.565 -12.075 ;
        RECT 596.875 -12.405 597.205 -12.075 ;
        RECT 595.515 -12.405 595.845 -12.075 ;
        RECT 594.155 -12.405 594.485 -12.075 ;
        RECT 592.795 -12.405 593.125 -12.075 ;
        RECT 591.435 -12.405 591.765 -12.075 ;
        RECT 590.075 -12.405 590.405 -12.075 ;
        RECT 588.715 -12.405 589.045 -12.075 ;
        RECT 587.355 -12.405 587.685 -12.075 ;
        RECT 585.995 -12.405 586.325 -12.075 ;
        RECT 584.635 -12.405 584.965 -12.075 ;
        RECT 583.275 -12.405 583.605 -12.075 ;
        RECT 581.915 -12.405 582.245 -12.075 ;
        RECT 580.555 -12.405 580.885 -12.075 ;
        RECT 579.195 -12.405 579.525 -12.075 ;
        RECT 577.835 -12.405 578.165 -12.075 ;
        RECT 576.475 -12.405 576.805 -12.075 ;
        RECT 575.115 -12.405 575.445 -12.075 ;
        RECT 573.755 -12.405 574.085 -12.075 ;
        RECT 572.395 -12.405 572.725 -12.075 ;
        RECT 571.035 -12.405 571.365 -12.075 ;
        RECT 569.675 -12.405 570.005 -12.075 ;
        RECT 568.315 -12.405 568.645 -12.075 ;
        RECT 566.955 -12.405 567.285 -12.075 ;
        RECT 565.595 -12.405 565.925 -12.075 ;
        RECT 564.235 -12.405 564.565 -12.075 ;
        RECT 562.875 -12.405 563.205 -12.075 ;
        RECT 561.515 -12.405 561.845 -12.075 ;
        RECT 560.155 -12.405 560.485 -12.075 ;
        RECT 558.795 -12.405 559.125 -12.075 ;
        RECT 557.435 -12.405 557.765 -12.075 ;
        RECT 556.075 -12.405 556.405 -12.075 ;
        RECT 554.715 -12.405 555.045 -12.075 ;
        RECT 553.355 -12.405 553.685 -12.075 ;
        RECT 551.995 -12.405 552.325 -12.075 ;
        RECT 550.635 -12.405 550.965 -12.075 ;
        RECT 549.275 -12.405 549.605 -12.075 ;
        RECT 547.915 -12.405 548.245 -12.075 ;
        RECT 546.555 -12.405 546.885 -12.075 ;
        RECT 545.195 -12.405 545.525 -12.075 ;
        RECT 543.835 -12.405 544.165 -12.075 ;
        RECT 542.475 -12.405 542.805 -12.075 ;
        RECT 541.115 -12.405 541.445 -12.075 ;
        RECT 539.755 -12.405 540.085 -12.075 ;
        RECT 538.395 -12.405 538.725 -12.075 ;
        RECT 537.035 -12.405 537.365 -12.075 ;
        RECT 535.675 -12.405 536.005 -12.075 ;
        RECT 534.315 -12.405 534.645 -12.075 ;
        RECT 532.955 -12.405 533.285 -12.075 ;
        RECT 531.595 -12.405 531.925 -12.075 ;
        RECT 530.235 -12.405 530.565 -12.075 ;
        RECT 528.875 -12.405 529.205 -12.075 ;
        RECT 527.515 -12.405 527.845 -12.075 ;
        RECT 526.155 -12.405 526.485 -12.075 ;
        RECT 524.795 -12.405 525.125 -12.075 ;
        RECT 523.435 -12.405 523.765 -12.075 ;
        RECT 522.075 -12.405 522.405 -12.075 ;
        RECT 520.715 -12.405 521.045 -12.075 ;
        RECT 519.355 -12.405 519.685 -12.075 ;
        RECT 517.995 -12.405 518.325 -12.075 ;
        RECT 516.635 -12.405 516.965 -12.075 ;
        RECT 515.275 -12.405 515.605 -12.075 ;
        RECT 513.915 -12.405 514.245 -12.075 ;
        RECT 512.555 -12.405 512.885 -12.075 ;
        RECT 511.195 -12.405 511.525 -12.075 ;
        RECT 509.835 -12.405 510.165 -12.075 ;
        RECT 508.475 -12.405 508.805 -12.075 ;
        RECT 507.115 -12.405 507.445 -12.075 ;
        RECT 505.755 -12.405 506.085 -12.075 ;
        RECT 504.395 -12.405 504.725 -12.075 ;
        RECT 503.035 -12.405 503.365 -12.075 ;
        RECT 501.675 -12.405 502.005 -12.075 ;
        RECT 500.315 -12.405 500.645 -12.075 ;
        RECT 498.955 -12.405 499.285 -12.075 ;
        RECT 497.595 -12.405 497.925 -12.075 ;
        RECT 496.235 -12.405 496.565 -12.075 ;
        RECT 494.875 -12.405 495.205 -12.075 ;
        RECT 493.515 -12.405 493.845 -12.075 ;
        RECT 492.155 -12.405 492.485 -12.075 ;
        RECT 490.795 -12.405 491.125 -12.075 ;
        RECT 489.435 -12.405 489.765 -12.075 ;
        RECT 488.075 -12.405 488.405 -12.075 ;
        RECT 486.715 -12.405 487.045 -12.075 ;
        RECT 485.355 -12.405 485.685 -12.075 ;
        RECT 483.995 -12.405 484.325 -12.075 ;
        RECT 482.635 -12.405 482.965 -12.075 ;
        RECT 481.275 -12.405 481.605 -12.075 ;
        RECT 479.915 -12.405 480.245 -12.075 ;
        RECT 478.555 -12.405 478.885 -12.075 ;
        RECT 477.195 -12.405 477.525 -12.075 ;
        RECT 475.835 -12.405 476.165 -12.075 ;
        RECT 474.475 -12.405 474.805 -12.075 ;
        RECT 473.115 -12.405 473.445 -12.075 ;
        RECT 471.755 -12.405 472.085 -12.075 ;
        RECT 470.395 -12.405 470.725 -12.075 ;
        RECT 469.035 -12.405 469.365 -12.075 ;
        RECT 467.675 -12.405 468.005 -12.075 ;
        RECT 466.315 -12.405 466.645 -12.075 ;
        RECT 464.955 -12.405 465.285 -12.075 ;
        RECT 463.595 -12.405 463.925 -12.075 ;
        RECT 462.235 -12.405 462.565 -12.075 ;
        RECT 460.875 -12.405 461.205 -12.075 ;
        RECT 459.515 -12.405 459.845 -12.075 ;
        RECT 458.155 -12.405 458.485 -12.075 ;
        RECT 456.795 -12.405 457.125 -12.075 ;
        RECT 455.435 -12.405 455.765 -12.075 ;
        RECT 454.075 -12.405 454.405 -12.075 ;
        RECT 452.715 -12.405 453.045 -12.075 ;
        RECT 451.355 -12.405 451.685 -12.075 ;
        RECT 449.995 -12.405 450.325 -12.075 ;
        RECT 448.635 -12.405 448.965 -12.075 ;
        RECT 447.275 -12.405 447.605 -12.075 ;
        RECT 445.915 -12.405 446.245 -12.075 ;
        RECT 444.555 -12.405 444.885 -12.075 ;
        RECT 443.195 -12.405 443.525 -12.075 ;
        RECT 441.835 -12.405 442.165 -12.075 ;
        RECT 440.475 -12.405 440.805 -12.075 ;
        RECT 439.115 -12.405 439.445 -12.075 ;
        RECT 437.755 -12.405 438.085 -12.075 ;
        RECT 436.395 -12.405 436.725 -12.075 ;
        RECT 435.035 -12.405 435.365 -12.075 ;
        RECT 433.675 -12.405 434.005 -12.075 ;
        RECT 432.315 -12.405 432.645 -12.075 ;
        RECT 430.955 -12.405 431.285 -12.075 ;
        RECT 429.595 -12.405 429.925 -12.075 ;
        RECT 428.235 -12.405 428.565 -12.075 ;
        RECT 426.875 -12.405 427.205 -12.075 ;
        RECT 425.515 -12.405 425.845 -12.075 ;
        RECT 424.155 -12.405 424.485 -12.075 ;
        RECT 422.795 -12.405 423.125 -12.075 ;
        RECT 421.435 -12.405 421.765 -12.075 ;
        RECT 420.075 -12.405 420.405 -12.075 ;
        RECT 418.715 -12.405 419.045 -12.075 ;
        RECT 417.355 -12.405 417.685 -12.075 ;
        RECT 415.995 -12.405 416.325 -12.075 ;
        RECT 414.635 -12.405 414.965 -12.075 ;
        RECT 413.275 -12.405 413.605 -12.075 ;
        RECT 411.915 -12.405 412.245 -12.075 ;
        RECT 410.555 -12.405 410.885 -12.075 ;
        RECT 409.195 -12.405 409.525 -12.075 ;
        RECT 407.835 -12.405 408.165 -12.075 ;
        RECT 406.475 -12.405 406.805 -12.075 ;
        RECT 405.115 -12.405 405.445 -12.075 ;
        RECT 403.755 -12.405 404.085 -12.075 ;
        RECT 402.395 -12.405 402.725 -12.075 ;
        RECT 401.035 -12.405 401.365 -12.075 ;
        RECT 399.675 -12.405 400.005 -12.075 ;
        RECT 398.315 -12.405 398.645 -12.075 ;
        RECT 396.955 -12.405 397.285 -12.075 ;
        RECT 395.595 -12.405 395.925 -12.075 ;
        RECT 394.235 -12.405 394.565 -12.075 ;
        RECT 392.875 -12.405 393.205 -12.075 ;
        RECT 391.515 -12.405 391.845 -12.075 ;
        RECT 390.155 -12.405 390.485 -12.075 ;
        RECT 388.795 -12.405 389.125 -12.075 ;
        RECT 387.435 -12.405 387.765 -12.075 ;
        RECT 386.075 -12.405 386.405 -12.075 ;
        RECT 384.715 -12.405 385.045 -12.075 ;
        RECT 383.355 -12.405 383.685 -12.075 ;
        RECT 381.995 -12.405 382.325 -12.075 ;
        RECT 380.635 -12.405 380.965 -12.075 ;
        RECT 379.275 -12.405 379.605 -12.075 ;
        RECT 377.915 -12.405 378.245 -12.075 ;
        RECT 376.555 -12.405 376.885 -12.075 ;
        RECT 375.195 -12.405 375.525 -12.075 ;
        RECT 373.835 -12.405 374.165 -12.075 ;
        RECT 372.475 -12.405 372.805 -12.075 ;
        RECT 371.115 -12.405 371.445 -12.075 ;
        RECT 369.755 -12.405 370.085 -12.075 ;
        RECT 368.395 -12.405 368.725 -12.075 ;
        RECT 367.035 -12.405 367.365 -12.075 ;
        RECT 365.675 -12.405 366.005 -12.075 ;
        RECT 364.315 -12.405 364.645 -12.075 ;
        RECT 362.955 -12.405 363.285 -12.075 ;
        RECT 361.595 -12.405 361.925 -12.075 ;
        RECT 360.235 -12.405 360.565 -12.075 ;
        RECT 358.875 -12.405 359.205 -12.075 ;
        RECT 357.515 -12.405 357.845 -12.075 ;
        RECT 356.155 -12.405 356.485 -12.075 ;
        RECT 354.795 -12.405 355.125 -12.075 ;
        RECT 353.435 -12.405 353.765 -12.075 ;
        RECT 352.075 -12.405 352.405 -12.075 ;
        RECT 350.715 -12.405 351.045 -12.075 ;
        RECT 349.355 -12.405 349.685 -12.075 ;
        RECT 347.995 -12.405 348.325 -12.075 ;
        RECT 346.635 -12.405 346.965 -12.075 ;
        RECT 345.275 -12.405 345.605 -12.075 ;
        RECT 343.915 -12.405 344.245 -12.075 ;
        RECT 342.555 -12.405 342.885 -12.075 ;
        RECT 341.195 -12.405 341.525 -12.075 ;
        RECT 339.835 -12.405 340.165 -12.075 ;
        RECT 338.475 -12.405 338.805 -12.075 ;
        RECT 337.115 -12.405 337.445 -12.075 ;
        RECT 335.755 -12.405 336.085 -12.075 ;
        RECT 334.395 -12.405 334.725 -12.075 ;
        RECT 333.035 -12.405 333.365 -12.075 ;
        RECT 331.675 -12.405 332.005 -12.075 ;
        RECT 330.315 -12.405 330.645 -12.075 ;
        RECT 328.955 -12.405 329.285 -12.075 ;
        RECT 327.595 -12.405 327.925 -12.075 ;
        RECT 326.235 -12.405 326.565 -12.075 ;
        RECT 324.875 -12.405 325.205 -12.075 ;
        RECT 323.515 -12.405 323.845 -12.075 ;
        RECT 322.155 -12.405 322.485 -12.075 ;
        RECT 320.795 -12.405 321.125 -12.075 ;
        RECT 319.435 -12.405 319.765 -12.075 ;
        RECT 318.075 -12.405 318.405 -12.075 ;
        RECT 316.715 -12.405 317.045 -12.075 ;
        RECT 315.355 -12.405 315.685 -12.075 ;
        RECT 313.995 -12.405 314.325 -12.075 ;
        RECT 312.635 -12.405 312.965 -12.075 ;
        RECT 311.275 -12.405 311.605 -12.075 ;
        RECT 309.915 -12.405 310.245 -12.075 ;
        RECT 308.555 -12.405 308.885 -12.075 ;
        RECT 307.195 -12.405 307.525 -12.075 ;
        RECT 305.835 -12.405 306.165 -12.075 ;
        RECT 304.475 -12.405 304.805 -12.075 ;
        RECT 303.115 -12.405 303.445 -12.075 ;
        RECT 301.755 -12.405 302.085 -12.075 ;
        RECT 300.395 -12.405 300.725 -12.075 ;
        RECT 299.035 -12.405 299.365 -12.075 ;
        RECT 297.675 -12.405 298.005 -12.075 ;
        RECT 296.315 -12.405 296.645 -12.075 ;
        RECT 294.955 -12.405 295.285 -12.075 ;
        RECT 293.595 -12.405 293.925 -12.075 ;
        RECT 292.235 -12.405 292.565 -12.075 ;
        RECT 290.875 -12.405 291.205 -12.075 ;
        RECT 289.515 -12.405 289.845 -12.075 ;
        RECT 288.155 -12.405 288.485 -12.075 ;
        RECT 286.795 -12.405 287.125 -12.075 ;
        RECT 285.435 -12.405 285.765 -12.075 ;
        RECT 284.075 -12.405 284.405 -12.075 ;
        RECT 282.715 -12.405 283.045 -12.075 ;
        RECT 281.355 -12.405 281.685 -12.075 ;
        RECT 279.995 -12.405 280.325 -12.075 ;
        RECT 278.635 -12.405 278.965 -12.075 ;
        RECT 277.275 -12.405 277.605 -12.075 ;
        RECT 275.915 -12.405 276.245 -12.075 ;
        RECT 274.555 -12.405 274.885 -12.075 ;
        RECT 273.195 -12.405 273.525 -12.075 ;
        RECT 271.835 -12.405 272.165 -12.075 ;
        RECT 270.475 -12.405 270.805 -12.075 ;
        RECT 269.115 -12.405 269.445 -12.075 ;
        RECT 267.755 -12.405 268.085 -12.075 ;
        RECT 266.395 -12.405 266.725 -12.075 ;
        RECT 265.035 -12.405 265.365 -12.075 ;
        RECT 263.675 -12.405 264.005 -12.075 ;
        RECT 262.315 -12.405 262.645 -12.075 ;
        RECT 260.955 -12.405 261.285 -12.075 ;
        RECT 259.595 -12.405 259.925 -12.075 ;
        RECT 258.235 -12.405 258.565 -12.075 ;
        RECT 256.875 -12.405 257.205 -12.075 ;
        RECT 255.515 -12.405 255.845 -12.075 ;
        RECT 254.155 -12.405 254.485 -12.075 ;
        RECT 252.795 -12.405 253.125 -12.075 ;
        RECT 251.435 -12.405 251.765 -12.075 ;
        RECT 250.075 -12.405 250.405 -12.075 ;
        RECT 248.715 -12.405 249.045 -12.075 ;
        RECT 247.355 -12.405 247.685 -12.075 ;
        RECT 245.995 -12.405 246.325 -12.075 ;
        RECT 244.635 -12.405 244.965 -12.075 ;
        RECT 243.275 -12.405 243.605 -12.075 ;
        RECT 241.915 -12.405 242.245 -12.075 ;
        RECT 240.555 -12.405 240.885 -12.075 ;
        RECT 239.195 -12.405 239.525 -12.075 ;
        RECT 237.835 -12.405 238.165 -12.075 ;
        RECT 236.475 -12.405 236.805 -12.075 ;
        RECT 235.115 -12.405 235.445 -12.075 ;
        RECT 233.755 -12.405 234.085 -12.075 ;
        RECT 232.395 -12.405 232.725 -12.075 ;
        RECT 231.035 -12.405 231.365 -12.075 ;
        RECT 229.675 -12.405 230.005 -12.075 ;
        RECT 228.315 -12.405 228.645 -12.075 ;
        RECT 226.955 -12.405 227.285 -12.075 ;
        RECT 225.595 -12.405 225.925 -12.075 ;
        RECT 224.235 -12.405 224.565 -12.075 ;
        RECT 222.875 -12.405 223.205 -12.075 ;
        RECT 221.515 -12.405 221.845 -12.075 ;
        RECT 220.155 -12.405 220.485 -12.075 ;
        RECT 218.795 -12.405 219.125 -12.075 ;
        RECT 217.435 -12.405 217.765 -12.075 ;
        RECT 216.075 -12.405 216.405 -12.075 ;
        RECT 214.715 -12.405 215.045 -12.075 ;
        RECT 213.355 -12.405 213.685 -12.075 ;
        RECT 211.995 -12.405 212.325 -12.075 ;
        RECT 210.635 -12.405 210.965 -12.075 ;
        RECT 209.275 -12.405 209.605 -12.075 ;
        RECT 207.915 -12.405 208.245 -12.075 ;
        RECT 206.555 -12.405 206.885 -12.075 ;
        RECT 205.195 -12.405 205.525 -12.075 ;
        RECT 203.835 -12.405 204.165 -12.075 ;
        RECT 202.475 -12.405 202.805 -12.075 ;
        RECT 201.115 -12.405 201.445 -12.075 ;
        RECT 199.755 -12.405 200.085 -12.075 ;
        RECT 198.395 -12.405 198.725 -12.075 ;
        RECT 197.035 -12.405 197.365 -12.075 ;
        RECT 195.675 -12.405 196.005 -12.075 ;
        RECT 194.315 -12.405 194.645 -12.075 ;
        RECT 192.955 -12.405 193.285 -12.075 ;
        RECT 191.595 -12.405 191.925 -12.075 ;
        RECT 190.235 -12.405 190.565 -12.075 ;
        RECT 188.875 -12.405 189.205 -12.075 ;
        RECT 187.515 -12.405 187.845 -12.075 ;
        RECT 186.155 -12.405 186.485 -12.075 ;
        RECT 184.795 -12.405 185.125 -12.075 ;
        RECT 183.435 -12.405 183.765 -12.075 ;
        RECT 182.075 -12.405 182.405 -12.075 ;
        RECT 180.715 -12.405 181.045 -12.075 ;
        RECT 179.355 -12.405 179.685 -12.075 ;
        RECT 177.995 -12.405 178.325 -12.075 ;
        RECT 176.635 -12.405 176.965 -12.075 ;
        RECT 175.275 -12.405 175.605 -12.075 ;
        RECT 173.915 -12.405 174.245 -12.075 ;
        RECT 172.555 -12.405 172.885 -12.075 ;
        RECT 171.195 -12.405 171.525 -12.075 ;
        RECT 169.835 -12.405 170.165 -12.075 ;
        RECT 168.475 -12.405 168.805 -12.075 ;
        RECT 167.115 -12.405 167.445 -12.075 ;
        RECT 165.755 -12.405 166.085 -12.075 ;
        RECT 164.395 -12.405 164.725 -12.075 ;
        RECT 163.035 -12.405 163.365 -12.075 ;
        RECT 161.675 -12.405 162.005 -12.075 ;
        RECT 160.315 -12.405 160.645 -12.075 ;
        RECT 158.955 -12.405 159.285 -12.075 ;
        RECT 157.595 -12.405 157.925 -12.075 ;
        RECT 156.235 -12.405 156.565 -12.075 ;
        RECT 154.875 -12.405 155.205 -12.075 ;
        RECT 153.515 -12.405 153.845 -12.075 ;
        RECT 152.155 -12.405 152.485 -12.075 ;
        RECT 150.795 -12.405 151.125 -12.075 ;
        RECT 149.435 -12.405 149.765 -12.075 ;
        RECT 148.075 -12.405 148.405 -12.075 ;
        RECT 146.715 -12.405 147.045 -12.075 ;
        RECT 145.355 -12.405 145.685 -12.075 ;
        RECT 143.995 -12.405 144.325 -12.075 ;
        RECT 142.635 -12.405 142.965 -12.075 ;
        RECT 141.275 -12.405 141.605 -12.075 ;
        RECT 139.915 -12.405 140.245 -12.075 ;
        RECT 138.555 -12.405 138.885 -12.075 ;
        RECT 137.195 -12.405 137.525 -12.075 ;
        RECT 135.835 -12.405 136.165 -12.075 ;
        RECT 134.475 -12.405 134.805 -12.075 ;
        RECT 133.115 -12.405 133.445 -12.075 ;
        RECT 131.755 -12.405 132.085 -12.075 ;
        RECT 130.395 -12.405 130.725 -12.075 ;
        RECT 129.035 -12.405 129.365 -12.075 ;
        RECT 127.675 -12.405 128.005 -12.075 ;
        RECT 126.315 -12.405 126.645 -12.075 ;
        RECT 124.955 -12.405 125.285 -12.075 ;
        RECT 123.595 -12.405 123.925 -12.075 ;
        RECT 122.235 -12.405 122.565 -12.075 ;
        RECT 120.875 -12.405 121.205 -12.075 ;
        RECT 119.515 -12.405 119.845 -12.075 ;
        RECT 118.155 -12.405 118.485 -12.075 ;
        RECT 116.795 -12.405 117.125 -12.075 ;
        RECT 115.435 -12.405 115.765 -12.075 ;
        RECT 114.075 -12.405 114.405 -12.075 ;
        RECT 112.715 -12.405 113.045 -12.075 ;
        RECT 111.355 -12.405 111.685 -12.075 ;
        RECT 109.995 -12.405 110.325 -12.075 ;
        RECT 108.635 -12.405 108.965 -12.075 ;
        RECT 107.275 -12.405 107.605 -12.075 ;
        RECT 105.915 -12.405 106.245 -12.075 ;
        RECT 104.555 -12.405 104.885 -12.075 ;
        RECT 103.195 -12.405 103.525 -12.075 ;
        RECT 101.835 -12.405 102.165 -12.075 ;
        RECT 100.475 -12.405 100.805 -12.075 ;
        RECT 99.115 -12.405 99.445 -12.075 ;
        RECT 97.755 -12.405 98.085 -12.075 ;
        RECT 96.395 -12.405 96.725 -12.075 ;
        RECT 95.035 -12.405 95.365 -12.075 ;
        RECT 93.675 -12.405 94.005 -12.075 ;
        RECT 92.315 -12.405 92.645 -12.075 ;
        RECT 90.955 -12.405 91.285 -12.075 ;
        RECT 89.595 -12.405 89.925 -12.075 ;
        RECT 88.235 -12.405 88.565 -12.075 ;
        RECT 86.875 -12.405 87.205 -12.075 ;
        RECT 85.515 -12.405 85.845 -12.075 ;
        RECT 84.155 -12.405 84.485 -12.075 ;
        RECT 82.795 -12.405 83.125 -12.075 ;
        RECT 81.435 -12.405 81.765 -12.075 ;
        RECT 80.075 -12.405 80.405 -12.075 ;
        RECT 78.715 -12.405 79.045 -12.075 ;
        RECT 77.355 -12.405 77.685 -12.075 ;
        RECT 75.995 -12.405 76.325 -12.075 ;
        RECT 74.635 -12.405 74.965 -12.075 ;
        RECT 73.275 -12.405 73.605 -12.075 ;
        RECT 71.915 -12.405 72.245 -12.075 ;
        RECT 70.555 -12.405 70.885 -12.075 ;
        RECT 69.195 -12.405 69.525 -12.075 ;
        RECT 67.835 -12.405 68.165 -12.075 ;
        RECT 66.475 -12.405 66.805 -12.075 ;
        RECT 65.115 -12.405 65.445 -12.075 ;
        RECT 63.755 -12.405 64.085 -12.075 ;
        RECT 62.395 -12.405 62.725 -12.075 ;
        RECT 61.035 -12.405 61.365 -12.075 ;
        RECT 59.675 -12.405 60.005 -12.075 ;
        RECT 58.315 -12.405 58.645 -12.075 ;
        RECT 56.955 -12.405 57.285 -12.075 ;
        RECT 55.595 -12.405 55.925 -12.075 ;
        RECT 54.235 -12.405 54.565 -12.075 ;
        RECT 52.875 -12.405 53.205 -12.075 ;
        RECT 51.515 -12.405 51.845 -12.075 ;
        RECT 50.155 -12.405 50.485 -12.075 ;
        RECT 48.795 -12.405 49.125 -12.075 ;
        RECT 47.435 -12.405 47.765 -12.075 ;
        RECT 46.075 -12.405 46.405 -12.075 ;
        RECT 44.715 -12.405 45.045 -12.075 ;
        RECT 43.355 -12.405 43.685 -12.075 ;
        RECT 41.995 -12.405 42.325 -12.075 ;
        RECT 40.635 -12.405 40.965 -12.075 ;
        RECT 39.275 -12.405 39.605 -12.075 ;
        RECT 37.915 -12.405 38.245 -12.075 ;
        RECT 36.555 -12.405 36.885 -12.075 ;
        RECT 35.195 -12.405 35.525 -12.075 ;
        RECT 33.835 -12.405 34.165 -12.075 ;
        RECT 32.475 -12.405 32.805 -12.075 ;
        RECT 31.115 -12.405 31.445 -12.075 ;
        RECT 29.755 -12.405 30.085 -12.075 ;
        RECT 28.395 -12.405 28.725 -12.075 ;
        RECT 27.035 -12.405 27.365 -12.075 ;
        RECT 25.675 -12.405 26.005 -12.075 ;
        RECT 24.315 -12.405 24.645 -12.075 ;
        RECT 22.955 -12.405 23.285 -12.075 ;
        RECT 21.595 -12.405 21.925 -12.075 ;
        RECT 20.235 -12.405 20.565 -12.075 ;
        RECT 18.875 -12.405 19.205 -12.075 ;
        RECT 17.515 -12.405 17.845 -12.075 ;
        RECT 16.155 -12.405 16.485 -12.075 ;
        RECT 14.795 -12.405 15.125 -12.075 ;
        RECT 13.435 -12.405 13.765 -12.075 ;
        RECT 12.075 -12.405 12.405 -12.075 ;
        RECT 10.715 -12.405 11.045 -12.075 ;
        RECT 9.355 -12.405 9.685 -12.075 ;
        RECT 7.995 -12.405 8.325 -12.075 ;
        RECT 6.635 -12.405 6.965 -12.075 ;
        RECT 5.275 -12.405 5.605 -12.075 ;
        RECT 3.915 -12.405 4.245 -12.075 ;
        RECT 2.555 -12.405 2.885 -12.075 ;
        RECT 1.195 -12.405 1.525 -12.075 ;
        RECT -0.165 -12.405 0.165 -12.075 ;
        RECT -1.525 -12.405 -1.195 -12.075 ;
        RECT 954.555 -12.405 954.885 -12.075 ;
        RECT 678.475 -12.4 954.885 -12.08 ;
        RECT 953.195 -12.405 953.525 -12.075 ;
        RECT 951.835 -12.405 952.165 -12.075 ;
        RECT 950.475 -12.405 950.805 -12.075 ;
        RECT 949.115 -12.405 949.445 -12.075 ;
        RECT 947.755 -12.405 948.085 -12.075 ;
        RECT 946.395 -12.405 946.725 -12.075 ;
        RECT 945.035 -12.405 945.365 -12.075 ;
        RECT 943.675 -12.405 944.005 -12.075 ;
        RECT 942.315 -12.405 942.645 -12.075 ;
        RECT 940.955 -12.405 941.285 -12.075 ;
        RECT 939.595 -12.405 939.925 -12.075 ;
        RECT 938.235 -12.405 938.565 -12.075 ;
        RECT 936.875 -12.405 937.205 -12.075 ;
        RECT 935.515 -12.405 935.845 -12.075 ;
        RECT 934.155 -12.405 934.485 -12.075 ;
        RECT 932.795 -12.405 933.125 -12.075 ;
        RECT 931.435 -12.405 931.765 -12.075 ;
        RECT 930.075 -12.405 930.405 -12.075 ;
        RECT 928.715 -12.405 929.045 -12.075 ;
        RECT 927.355 -12.405 927.685 -12.075 ;
        RECT 925.995 -12.405 926.325 -12.075 ;
        RECT 924.635 -12.405 924.965 -12.075 ;
        RECT 923.275 -12.405 923.605 -12.075 ;
        RECT 921.915 -12.405 922.245 -12.075 ;
        RECT 920.555 -12.405 920.885 -12.075 ;
        RECT 919.195 -12.405 919.525 -12.075 ;
        RECT 917.835 -12.405 918.165 -12.075 ;
        RECT 916.475 -12.405 916.805 -12.075 ;
        RECT 915.115 -12.405 915.445 -12.075 ;
        RECT 913.755 -12.405 914.085 -12.075 ;
        RECT 912.395 -12.405 912.725 -12.075 ;
        RECT 911.035 -12.405 911.365 -12.075 ;
        RECT 909.675 -12.405 910.005 -12.075 ;
        RECT 908.315 -12.405 908.645 -12.075 ;
        RECT 906.955 -12.405 907.285 -12.075 ;
        RECT 905.595 -12.405 905.925 -12.075 ;
        RECT 904.235 -12.405 904.565 -12.075 ;
        RECT 902.875 -12.405 903.205 -12.075 ;
        RECT 901.515 -12.405 901.845 -12.075 ;
        RECT 900.155 -12.405 900.485 -12.075 ;
        RECT 898.795 -12.405 899.125 -12.075 ;
        RECT 897.435 -12.405 897.765 -12.075 ;
        RECT 896.075 -12.405 896.405 -12.075 ;
        RECT 894.715 -12.405 895.045 -12.075 ;
        RECT 893.355 -12.405 893.685 -12.075 ;
        RECT 891.995 -12.405 892.325 -12.075 ;
        RECT 890.635 -12.405 890.965 -12.075 ;
        RECT 889.275 -12.405 889.605 -12.075 ;
        RECT 887.915 -12.405 888.245 -12.075 ;
        RECT 886.555 -12.405 886.885 -12.075 ;
        RECT 885.195 -12.405 885.525 -12.075 ;
        RECT 883.835 -12.405 884.165 -12.075 ;
        RECT 882.475 -12.405 882.805 -12.075 ;
        RECT 881.115 -12.405 881.445 -12.075 ;
        RECT 879.755 -12.405 880.085 -12.075 ;
        RECT 878.395 -12.405 878.725 -12.075 ;
        RECT 877.035 -12.405 877.365 -12.075 ;
        RECT 875.675 -12.405 876.005 -12.075 ;
        RECT 874.315 -12.405 874.645 -12.075 ;
        RECT 872.955 -12.405 873.285 -12.075 ;
        RECT 871.595 -12.405 871.925 -12.075 ;
        RECT 870.235 -12.405 870.565 -12.075 ;
        RECT 868.875 -12.405 869.205 -12.075 ;
        RECT 867.515 -12.405 867.845 -12.075 ;
        RECT 866.155 -12.405 866.485 -12.075 ;
        RECT 864.795 -12.405 865.125 -12.075 ;
        RECT 863.435 -12.405 863.765 -12.075 ;
        RECT 862.075 -12.405 862.405 -12.075 ;
        RECT 860.715 -12.405 861.045 -12.075 ;
        RECT 859.355 -12.405 859.685 -12.075 ;
        RECT 857.995 -12.405 858.325 -12.075 ;
        RECT 856.635 -12.405 856.965 -12.075 ;
        RECT 855.275 -12.405 855.605 -12.075 ;
        RECT 853.915 -12.405 854.245 -12.075 ;
        RECT 852.555 -12.405 852.885 -12.075 ;
        RECT 851.195 -12.405 851.525 -12.075 ;
        RECT 849.835 -12.405 850.165 -12.075 ;
        RECT 848.475 -12.405 848.805 -12.075 ;
        RECT 847.115 -12.405 847.445 -12.075 ;
        RECT 845.755 -12.405 846.085 -12.075 ;
        RECT 844.395 -12.405 844.725 -12.075 ;
        RECT 843.035 -12.405 843.365 -12.075 ;
        RECT 841.675 -12.405 842.005 -12.075 ;
        RECT 840.315 -12.405 840.645 -12.075 ;
        RECT 838.955 -12.405 839.285 -12.075 ;
        RECT 837.595 -12.405 837.925 -12.075 ;
        RECT 836.235 -12.405 836.565 -12.075 ;
        RECT 834.875 -12.405 835.205 -12.075 ;
        RECT 833.515 -12.405 833.845 -12.075 ;
        RECT 832.155 -12.405 832.485 -12.075 ;
        RECT 830.795 -12.405 831.125 -12.075 ;
        RECT 829.435 -12.405 829.765 -12.075 ;
        RECT 828.075 -12.405 828.405 -12.075 ;
        RECT 826.715 -12.405 827.045 -12.075 ;
        RECT 825.355 -12.405 825.685 -12.075 ;
        RECT 823.995 -12.405 824.325 -12.075 ;
        RECT 822.635 -12.405 822.965 -12.075 ;
        RECT 821.275 -12.405 821.605 -12.075 ;
        RECT 819.915 -12.405 820.245 -12.075 ;
        RECT 818.555 -12.405 818.885 -12.075 ;
        RECT 817.195 -12.405 817.525 -12.075 ;
        RECT 815.835 -12.405 816.165 -12.075 ;
        RECT 814.475 -12.405 814.805 -12.075 ;
        RECT 813.115 -12.405 813.445 -12.075 ;
        RECT 811.755 -12.405 812.085 -12.075 ;
        RECT 810.395 -12.405 810.725 -12.075 ;
        RECT 809.035 -12.405 809.365 -12.075 ;
        RECT 807.675 -12.405 808.005 -12.075 ;
        RECT 806.315 -12.405 806.645 -12.075 ;
        RECT 804.955 -12.405 805.285 -12.075 ;
        RECT 803.595 -12.405 803.925 -12.075 ;
        RECT 802.235 -12.405 802.565 -12.075 ;
        RECT 800.875 -12.405 801.205 -12.075 ;
        RECT 799.515 -12.405 799.845 -12.075 ;
        RECT 798.155 -12.405 798.485 -12.075 ;
        RECT 796.795 -12.405 797.125 -12.075 ;
        RECT 795.435 -12.405 795.765 -12.075 ;
        RECT 794.075 -12.405 794.405 -12.075 ;
        RECT 792.715 -12.405 793.045 -12.075 ;
        RECT 791.355 -12.405 791.685 -12.075 ;
        RECT 789.995 -12.405 790.325 -12.075 ;
        RECT 788.635 -12.405 788.965 -12.075 ;
        RECT 787.275 -12.405 787.605 -12.075 ;
        RECT 785.915 -12.405 786.245 -12.075 ;
        RECT 784.555 -12.405 784.885 -12.075 ;
        RECT 783.195 -12.405 783.525 -12.075 ;
        RECT 781.835 -12.405 782.165 -12.075 ;
        RECT 780.475 -12.405 780.805 -12.075 ;
        RECT 779.115 -12.405 779.445 -12.075 ;
        RECT 777.755 -12.405 778.085 -12.075 ;
        RECT 776.395 -12.405 776.725 -12.075 ;
        RECT 775.035 -12.405 775.365 -12.075 ;
        RECT 773.675 -12.405 774.005 -12.075 ;
        RECT 772.315 -12.405 772.645 -12.075 ;
        RECT 770.955 -12.405 771.285 -12.075 ;
        RECT 769.595 -12.405 769.925 -12.075 ;
        RECT 768.235 -12.405 768.565 -12.075 ;
        RECT 766.875 -12.405 767.205 -12.075 ;
        RECT 765.515 -12.405 765.845 -12.075 ;
        RECT 764.155 -12.405 764.485 -12.075 ;
        RECT 762.795 -12.405 763.125 -12.075 ;
        RECT 761.435 -12.405 761.765 -12.075 ;
        RECT 760.075 -12.405 760.405 -12.075 ;
        RECT 758.715 -12.405 759.045 -12.075 ;
        RECT 757.355 -12.405 757.685 -12.075 ;
        RECT 755.995 -12.405 756.325 -12.075 ;
        RECT 754.635 -12.405 754.965 -12.075 ;
        RECT 753.275 -12.405 753.605 -12.075 ;
        RECT 751.915 -12.405 752.245 -12.075 ;
        RECT 750.555 -12.405 750.885 -12.075 ;
        RECT 749.195 -12.405 749.525 -12.075 ;
        RECT 747.835 -12.405 748.165 -12.075 ;
        RECT 746.475 -12.405 746.805 -12.075 ;
        RECT 745.115 -12.405 745.445 -12.075 ;
        RECT 743.755 -12.405 744.085 -12.075 ;
        RECT 742.395 -12.405 742.725 -12.075 ;
        RECT 741.035 -12.405 741.365 -12.075 ;
        RECT 739.675 -12.405 740.005 -12.075 ;
        RECT 738.315 -12.405 738.645 -12.075 ;
        RECT 736.955 -12.405 737.285 -12.075 ;
        RECT 735.595 -12.405 735.925 -12.075 ;
        RECT 734.235 -12.405 734.565 -12.075 ;
        RECT 732.875 -12.405 733.205 -12.075 ;
        RECT 731.515 -12.405 731.845 -12.075 ;
        RECT 730.155 -12.405 730.485 -12.075 ;
        RECT 728.795 -12.405 729.125 -12.075 ;
        RECT 727.435 -12.405 727.765 -12.075 ;
        RECT 726.075 -12.405 726.405 -12.075 ;
        RECT 724.715 -12.405 725.045 -12.075 ;
        RECT 723.355 -12.405 723.685 -12.075 ;
        RECT 721.995 -12.405 722.325 -12.075 ;
        RECT 720.635 -12.405 720.965 -12.075 ;
        RECT 719.275 -12.405 719.605 -12.075 ;
        RECT 717.915 -12.405 718.245 -12.075 ;
        RECT 716.555 -12.405 716.885 -12.075 ;
        RECT 715.195 -12.405 715.525 -12.075 ;
        RECT 713.835 -12.405 714.165 -12.075 ;
        RECT 712.475 -12.405 712.805 -12.075 ;
        RECT 711.115 -12.405 711.445 -12.075 ;
        RECT 709.755 -12.405 710.085 -12.075 ;
        RECT 708.395 -12.405 708.725 -12.075 ;
        RECT 707.035 -12.405 707.365 -12.075 ;
        RECT 705.675 -12.405 706.005 -12.075 ;
        RECT 704.315 -12.405 704.645 -12.075 ;
        RECT 702.955 -12.405 703.285 -12.075 ;
        RECT 701.595 -12.405 701.925 -12.075 ;
        RECT 700.235 -12.405 700.565 -12.075 ;
        RECT 698.875 -12.405 699.205 -12.075 ;
        RECT 697.515 -12.405 697.845 -12.075 ;
        RECT 696.155 -12.405 696.485 -12.075 ;
        RECT 694.795 -12.405 695.125 -12.075 ;
        RECT 693.435 -12.405 693.765 -12.075 ;
        RECT 692.075 -12.405 692.405 -12.075 ;
        RECT 690.715 -12.405 691.045 -12.075 ;
        RECT 689.355 -12.405 689.685 -12.075 ;
        RECT 687.995 -12.405 688.325 -12.075 ;
        RECT 686.635 -12.405 686.965 -12.075 ;
        RECT 685.275 -12.405 685.605 -12.075 ;
        RECT 683.915 -12.405 684.245 -12.075 ;
        RECT 682.555 -12.405 682.885 -12.075 ;
        RECT 681.195 -12.405 681.525 -12.075 ;
        RECT 679.835 -12.405 680.165 -12.075 ;
        RECT 678.475 -12.405 678.805 -12.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 645.835 -13.765 646.165 -13.435 ;
        RECT 644.475 -13.765 644.805 -13.435 ;
        RECT 643.115 -13.765 643.445 -13.435 ;
        RECT 641.755 -13.765 642.085 -13.435 ;
        RECT 640.395 -13.765 640.725 -13.435 ;
        RECT 639.035 -13.765 639.365 -13.435 ;
        RECT 637.675 -13.765 638.005 -13.435 ;
        RECT 636.315 -13.765 636.645 -13.435 ;
        RECT 634.955 -13.765 635.285 -13.435 ;
        RECT 633.595 -13.765 633.925 -13.435 ;
        RECT 632.235 -13.765 632.565 -13.435 ;
        RECT 630.875 -13.765 631.205 -13.435 ;
        RECT 629.515 -13.765 629.845 -13.435 ;
        RECT 628.155 -13.765 628.485 -13.435 ;
        RECT 626.795 -13.765 627.125 -13.435 ;
        RECT 625.435 -13.765 625.765 -13.435 ;
        RECT 624.075 -13.765 624.405 -13.435 ;
        RECT 622.715 -13.765 623.045 -13.435 ;
        RECT 621.355 -13.765 621.685 -13.435 ;
        RECT 619.995 -13.765 620.325 -13.435 ;
        RECT 618.635 -13.765 618.965 -13.435 ;
        RECT 617.275 -13.765 617.605 -13.435 ;
        RECT 615.915 -13.765 616.245 -13.435 ;
        RECT 614.555 -13.765 614.885 -13.435 ;
        RECT 613.195 -13.765 613.525 -13.435 ;
        RECT 611.835 -13.765 612.165 -13.435 ;
        RECT 610.475 -13.765 610.805 -13.435 ;
        RECT 609.115 -13.765 609.445 -13.435 ;
        RECT 607.755 -13.765 608.085 -13.435 ;
        RECT 606.395 -13.765 606.725 -13.435 ;
        RECT 605.035 -13.765 605.365 -13.435 ;
        RECT 603.675 -13.765 604.005 -13.435 ;
        RECT 602.315 -13.765 602.645 -13.435 ;
        RECT 600.955 -13.765 601.285 -13.435 ;
        RECT 599.595 -13.765 599.925 -13.435 ;
        RECT 598.235 -13.765 598.565 -13.435 ;
        RECT 596.875 -13.765 597.205 -13.435 ;
        RECT 595.515 -13.765 595.845 -13.435 ;
        RECT 594.155 -13.765 594.485 -13.435 ;
        RECT 592.795 -13.765 593.125 -13.435 ;
        RECT 591.435 -13.765 591.765 -13.435 ;
        RECT 590.075 -13.765 590.405 -13.435 ;
        RECT 588.715 -13.765 589.045 -13.435 ;
        RECT 587.355 -13.765 587.685 -13.435 ;
        RECT 585.995 -13.765 586.325 -13.435 ;
        RECT 584.635 -13.765 584.965 -13.435 ;
        RECT 583.275 -13.765 583.605 -13.435 ;
        RECT 581.915 -13.765 582.245 -13.435 ;
        RECT 580.555 -13.765 580.885 -13.435 ;
        RECT 579.195 -13.765 579.525 -13.435 ;
        RECT 577.835 -13.765 578.165 -13.435 ;
        RECT 576.475 -13.765 576.805 -13.435 ;
        RECT 575.115 -13.765 575.445 -13.435 ;
        RECT 573.755 -13.765 574.085 -13.435 ;
        RECT 572.395 -13.765 572.725 -13.435 ;
        RECT 571.035 -13.765 571.365 -13.435 ;
        RECT 569.675 -13.765 570.005 -13.435 ;
        RECT 568.315 -13.765 568.645 -13.435 ;
        RECT 566.955 -13.765 567.285 -13.435 ;
        RECT 565.595 -13.765 565.925 -13.435 ;
        RECT 564.235 -13.765 564.565 -13.435 ;
        RECT 562.875 -13.765 563.205 -13.435 ;
        RECT 561.515 -13.765 561.845 -13.435 ;
        RECT 560.155 -13.765 560.485 -13.435 ;
        RECT 558.795 -13.765 559.125 -13.435 ;
        RECT 557.435 -13.765 557.765 -13.435 ;
        RECT 556.075 -13.765 556.405 -13.435 ;
        RECT 554.715 -13.765 555.045 -13.435 ;
        RECT 553.355 -13.765 553.685 -13.435 ;
        RECT 551.995 -13.765 552.325 -13.435 ;
        RECT 550.635 -13.765 550.965 -13.435 ;
        RECT 549.275 -13.765 549.605 -13.435 ;
        RECT 547.915 -13.765 548.245 -13.435 ;
        RECT 546.555 -13.765 546.885 -13.435 ;
        RECT 545.195 -13.765 545.525 -13.435 ;
        RECT 543.835 -13.765 544.165 -13.435 ;
        RECT 542.475 -13.765 542.805 -13.435 ;
        RECT 541.115 -13.765 541.445 -13.435 ;
        RECT 539.755 -13.765 540.085 -13.435 ;
        RECT 538.395 -13.765 538.725 -13.435 ;
        RECT 537.035 -13.765 537.365 -13.435 ;
        RECT 535.675 -13.765 536.005 -13.435 ;
        RECT 534.315 -13.765 534.645 -13.435 ;
        RECT 532.955 -13.765 533.285 -13.435 ;
        RECT 531.595 -13.765 531.925 -13.435 ;
        RECT 530.235 -13.765 530.565 -13.435 ;
        RECT 528.875 -13.765 529.205 -13.435 ;
        RECT 527.515 -13.765 527.845 -13.435 ;
        RECT 526.155 -13.765 526.485 -13.435 ;
        RECT 524.795 -13.765 525.125 -13.435 ;
        RECT 523.435 -13.765 523.765 -13.435 ;
        RECT 522.075 -13.765 522.405 -13.435 ;
        RECT 520.715 -13.765 521.045 -13.435 ;
        RECT 519.355 -13.765 519.685 -13.435 ;
        RECT 517.995 -13.765 518.325 -13.435 ;
        RECT 516.635 -13.765 516.965 -13.435 ;
        RECT 515.275 -13.765 515.605 -13.435 ;
        RECT 513.915 -13.765 514.245 -13.435 ;
        RECT 512.555 -13.765 512.885 -13.435 ;
        RECT 511.195 -13.765 511.525 -13.435 ;
        RECT 509.835 -13.765 510.165 -13.435 ;
        RECT 508.475 -13.765 508.805 -13.435 ;
        RECT 507.115 -13.765 507.445 -13.435 ;
        RECT 505.755 -13.765 506.085 -13.435 ;
        RECT 504.395 -13.765 504.725 -13.435 ;
        RECT 503.035 -13.765 503.365 -13.435 ;
        RECT 501.675 -13.765 502.005 -13.435 ;
        RECT 500.315 -13.765 500.645 -13.435 ;
        RECT 498.955 -13.765 499.285 -13.435 ;
        RECT 497.595 -13.765 497.925 -13.435 ;
        RECT 496.235 -13.765 496.565 -13.435 ;
        RECT 494.875 -13.765 495.205 -13.435 ;
        RECT 493.515 -13.765 493.845 -13.435 ;
        RECT 492.155 -13.765 492.485 -13.435 ;
        RECT 490.795 -13.765 491.125 -13.435 ;
        RECT 489.435 -13.765 489.765 -13.435 ;
        RECT 488.075 -13.765 488.405 -13.435 ;
        RECT 486.715 -13.765 487.045 -13.435 ;
        RECT 485.355 -13.765 485.685 -13.435 ;
        RECT 483.995 -13.765 484.325 -13.435 ;
        RECT 482.635 -13.765 482.965 -13.435 ;
        RECT 481.275 -13.765 481.605 -13.435 ;
        RECT 479.915 -13.765 480.245 -13.435 ;
        RECT 478.555 -13.765 478.885 -13.435 ;
        RECT 477.195 -13.765 477.525 -13.435 ;
        RECT 475.835 -13.765 476.165 -13.435 ;
        RECT 474.475 -13.765 474.805 -13.435 ;
        RECT 473.115 -13.765 473.445 -13.435 ;
        RECT 471.755 -13.765 472.085 -13.435 ;
        RECT 470.395 -13.765 470.725 -13.435 ;
        RECT 469.035 -13.765 469.365 -13.435 ;
        RECT 467.675 -13.765 468.005 -13.435 ;
        RECT 466.315 -13.765 466.645 -13.435 ;
        RECT 464.955 -13.765 465.285 -13.435 ;
        RECT 463.595 -13.765 463.925 -13.435 ;
        RECT 462.235 -13.765 462.565 -13.435 ;
        RECT 460.875 -13.765 461.205 -13.435 ;
        RECT 459.515 -13.765 459.845 -13.435 ;
        RECT 458.155 -13.765 458.485 -13.435 ;
        RECT 456.795 -13.765 457.125 -13.435 ;
        RECT 455.435 -13.765 455.765 -13.435 ;
        RECT 454.075 -13.765 454.405 -13.435 ;
        RECT 452.715 -13.765 453.045 -13.435 ;
        RECT 451.355 -13.765 451.685 -13.435 ;
        RECT 449.995 -13.765 450.325 -13.435 ;
        RECT 448.635 -13.765 448.965 -13.435 ;
        RECT 447.275 -13.765 447.605 -13.435 ;
        RECT 445.915 -13.765 446.245 -13.435 ;
        RECT 444.555 -13.765 444.885 -13.435 ;
        RECT 443.195 -13.765 443.525 -13.435 ;
        RECT 441.835 -13.765 442.165 -13.435 ;
        RECT 440.475 -13.765 440.805 -13.435 ;
        RECT 439.115 -13.765 439.445 -13.435 ;
        RECT 437.755 -13.765 438.085 -13.435 ;
        RECT 436.395 -13.765 436.725 -13.435 ;
        RECT 435.035 -13.765 435.365 -13.435 ;
        RECT 433.675 -13.765 434.005 -13.435 ;
        RECT 432.315 -13.765 432.645 -13.435 ;
        RECT 430.955 -13.765 431.285 -13.435 ;
        RECT 429.595 -13.765 429.925 -13.435 ;
        RECT 428.235 -13.765 428.565 -13.435 ;
        RECT 426.875 -13.765 427.205 -13.435 ;
        RECT 425.515 -13.765 425.845 -13.435 ;
        RECT 424.155 -13.765 424.485 -13.435 ;
        RECT 422.795 -13.765 423.125 -13.435 ;
        RECT 421.435 -13.765 421.765 -13.435 ;
        RECT 420.075 -13.765 420.405 -13.435 ;
        RECT 418.715 -13.765 419.045 -13.435 ;
        RECT 417.355 -13.765 417.685 -13.435 ;
        RECT 415.995 -13.765 416.325 -13.435 ;
        RECT 414.635 -13.765 414.965 -13.435 ;
        RECT 413.275 -13.765 413.605 -13.435 ;
        RECT 411.915 -13.765 412.245 -13.435 ;
        RECT 410.555 -13.765 410.885 -13.435 ;
        RECT 409.195 -13.765 409.525 -13.435 ;
        RECT 407.835 -13.765 408.165 -13.435 ;
        RECT 406.475 -13.765 406.805 -13.435 ;
        RECT 405.115 -13.765 405.445 -13.435 ;
        RECT 403.755 -13.765 404.085 -13.435 ;
        RECT 402.395 -13.765 402.725 -13.435 ;
        RECT 401.035 -13.765 401.365 -13.435 ;
        RECT 399.675 -13.765 400.005 -13.435 ;
        RECT 398.315 -13.765 398.645 -13.435 ;
        RECT 396.955 -13.765 397.285 -13.435 ;
        RECT 395.595 -13.765 395.925 -13.435 ;
        RECT 394.235 -13.765 394.565 -13.435 ;
        RECT 392.875 -13.765 393.205 -13.435 ;
        RECT 391.515 -13.765 391.845 -13.435 ;
        RECT 390.155 -13.765 390.485 -13.435 ;
        RECT 388.795 -13.765 389.125 -13.435 ;
        RECT 387.435 -13.765 387.765 -13.435 ;
        RECT 386.075 -13.765 386.405 -13.435 ;
        RECT 384.715 -13.765 385.045 -13.435 ;
        RECT 383.355 -13.765 383.685 -13.435 ;
        RECT 381.995 -13.765 382.325 -13.435 ;
        RECT 380.635 -13.765 380.965 -13.435 ;
        RECT 379.275 -13.765 379.605 -13.435 ;
        RECT 377.915 -13.765 378.245 -13.435 ;
        RECT 376.555 -13.765 376.885 -13.435 ;
        RECT 375.195 -13.765 375.525 -13.435 ;
        RECT 373.835 -13.765 374.165 -13.435 ;
        RECT 372.475 -13.765 372.805 -13.435 ;
        RECT 371.115 -13.765 371.445 -13.435 ;
        RECT 369.755 -13.765 370.085 -13.435 ;
        RECT 368.395 -13.765 368.725 -13.435 ;
        RECT 367.035 -13.765 367.365 -13.435 ;
        RECT 365.675 -13.765 366.005 -13.435 ;
        RECT 364.315 -13.765 364.645 -13.435 ;
        RECT 362.955 -13.765 363.285 -13.435 ;
        RECT 361.595 -13.765 361.925 -13.435 ;
        RECT 360.235 -13.765 360.565 -13.435 ;
        RECT 358.875 -13.765 359.205 -13.435 ;
        RECT 357.515 -13.765 357.845 -13.435 ;
        RECT 356.155 -13.765 356.485 -13.435 ;
        RECT 354.795 -13.765 355.125 -13.435 ;
        RECT 353.435 -13.765 353.765 -13.435 ;
        RECT 352.075 -13.765 352.405 -13.435 ;
        RECT 350.715 -13.765 351.045 -13.435 ;
        RECT 349.355 -13.765 349.685 -13.435 ;
        RECT 347.995 -13.765 348.325 -13.435 ;
        RECT 346.635 -13.765 346.965 -13.435 ;
        RECT 345.275 -13.765 345.605 -13.435 ;
        RECT 343.915 -13.765 344.245 -13.435 ;
        RECT 342.555 -13.765 342.885 -13.435 ;
        RECT 341.195 -13.765 341.525 -13.435 ;
        RECT 339.835 -13.765 340.165 -13.435 ;
        RECT 338.475 -13.765 338.805 -13.435 ;
        RECT 337.115 -13.765 337.445 -13.435 ;
        RECT 335.755 -13.765 336.085 -13.435 ;
        RECT 334.395 -13.765 334.725 -13.435 ;
        RECT 333.035 -13.765 333.365 -13.435 ;
        RECT 331.675 -13.765 332.005 -13.435 ;
        RECT 330.315 -13.765 330.645 -13.435 ;
        RECT 328.955 -13.765 329.285 -13.435 ;
        RECT 327.595 -13.765 327.925 -13.435 ;
        RECT 326.235 -13.765 326.565 -13.435 ;
        RECT 324.875 -13.765 325.205 -13.435 ;
        RECT 323.515 -13.765 323.845 -13.435 ;
        RECT 322.155 -13.765 322.485 -13.435 ;
        RECT 320.795 -13.765 321.125 -13.435 ;
        RECT 319.435 -13.765 319.765 -13.435 ;
        RECT 318.075 -13.765 318.405 -13.435 ;
        RECT 316.715 -13.765 317.045 -13.435 ;
        RECT 315.355 -13.765 315.685 -13.435 ;
        RECT 313.995 -13.765 314.325 -13.435 ;
        RECT 312.635 -13.765 312.965 -13.435 ;
        RECT 311.275 -13.765 311.605 -13.435 ;
        RECT 309.915 -13.765 310.245 -13.435 ;
        RECT 308.555 -13.765 308.885 -13.435 ;
        RECT 307.195 -13.765 307.525 -13.435 ;
        RECT 305.835 -13.765 306.165 -13.435 ;
        RECT 304.475 -13.765 304.805 -13.435 ;
        RECT 303.115 -13.765 303.445 -13.435 ;
        RECT 301.755 -13.765 302.085 -13.435 ;
        RECT 300.395 -13.765 300.725 -13.435 ;
        RECT 299.035 -13.765 299.365 -13.435 ;
        RECT 297.675 -13.765 298.005 -13.435 ;
        RECT 296.315 -13.765 296.645 -13.435 ;
        RECT 294.955 -13.765 295.285 -13.435 ;
        RECT 293.595 -13.765 293.925 -13.435 ;
        RECT 292.235 -13.765 292.565 -13.435 ;
        RECT 290.875 -13.765 291.205 -13.435 ;
        RECT 289.515 -13.765 289.845 -13.435 ;
        RECT 288.155 -13.765 288.485 -13.435 ;
        RECT 286.795 -13.765 287.125 -13.435 ;
        RECT 285.435 -13.765 285.765 -13.435 ;
        RECT 284.075 -13.765 284.405 -13.435 ;
        RECT 282.715 -13.765 283.045 -13.435 ;
        RECT 281.355 -13.765 281.685 -13.435 ;
        RECT 279.995 -13.765 280.325 -13.435 ;
        RECT 278.635 -13.765 278.965 -13.435 ;
        RECT 277.275 -13.765 277.605 -13.435 ;
        RECT 275.915 -13.765 276.245 -13.435 ;
        RECT 274.555 -13.765 274.885 -13.435 ;
        RECT 273.195 -13.765 273.525 -13.435 ;
        RECT 271.835 -13.765 272.165 -13.435 ;
        RECT 270.475 -13.765 270.805 -13.435 ;
        RECT 269.115 -13.765 269.445 -13.435 ;
        RECT 267.755 -13.765 268.085 -13.435 ;
        RECT 266.395 -13.765 266.725 -13.435 ;
        RECT 265.035 -13.765 265.365 -13.435 ;
        RECT 263.675 -13.765 264.005 -13.435 ;
        RECT 262.315 -13.765 262.645 -13.435 ;
        RECT 260.955 -13.765 261.285 -13.435 ;
        RECT 259.595 -13.765 259.925 -13.435 ;
        RECT 258.235 -13.765 258.565 -13.435 ;
        RECT 256.875 -13.765 257.205 -13.435 ;
        RECT 255.515 -13.765 255.845 -13.435 ;
        RECT 254.155 -13.765 254.485 -13.435 ;
        RECT 252.795 -13.765 253.125 -13.435 ;
        RECT 251.435 -13.765 251.765 -13.435 ;
        RECT 250.075 -13.765 250.405 -13.435 ;
        RECT 248.715 -13.765 249.045 -13.435 ;
        RECT 247.355 -13.765 247.685 -13.435 ;
        RECT 245.995 -13.765 246.325 -13.435 ;
        RECT 244.635 -13.765 244.965 -13.435 ;
        RECT 243.275 -13.765 243.605 -13.435 ;
        RECT 241.915 -13.765 242.245 -13.435 ;
        RECT 240.555 -13.765 240.885 -13.435 ;
        RECT 239.195 -13.765 239.525 -13.435 ;
        RECT 237.835 -13.765 238.165 -13.435 ;
        RECT 236.475 -13.765 236.805 -13.435 ;
        RECT 235.115 -13.765 235.445 -13.435 ;
        RECT 233.755 -13.765 234.085 -13.435 ;
        RECT 232.395 -13.765 232.725 -13.435 ;
        RECT 231.035 -13.765 231.365 -13.435 ;
        RECT 229.675 -13.765 230.005 -13.435 ;
        RECT 228.315 -13.765 228.645 -13.435 ;
        RECT 226.955 -13.765 227.285 -13.435 ;
        RECT 225.595 -13.765 225.925 -13.435 ;
        RECT 224.235 -13.765 224.565 -13.435 ;
        RECT 222.875 -13.765 223.205 -13.435 ;
        RECT 221.515 -13.765 221.845 -13.435 ;
        RECT 220.155 -13.765 220.485 -13.435 ;
        RECT 218.795 -13.765 219.125 -13.435 ;
        RECT 217.435 -13.765 217.765 -13.435 ;
        RECT 216.075 -13.765 216.405 -13.435 ;
        RECT 214.715 -13.765 215.045 -13.435 ;
        RECT 213.355 -13.765 213.685 -13.435 ;
        RECT 211.995 -13.765 212.325 -13.435 ;
        RECT 210.635 -13.765 210.965 -13.435 ;
        RECT 209.275 -13.765 209.605 -13.435 ;
        RECT 207.915 -13.765 208.245 -13.435 ;
        RECT 206.555 -13.765 206.885 -13.435 ;
        RECT 205.195 -13.765 205.525 -13.435 ;
        RECT 203.835 -13.765 204.165 -13.435 ;
        RECT 202.475 -13.765 202.805 -13.435 ;
        RECT 201.115 -13.765 201.445 -13.435 ;
        RECT 199.755 -13.765 200.085 -13.435 ;
        RECT 198.395 -13.765 198.725 -13.435 ;
        RECT 197.035 -13.765 197.365 -13.435 ;
        RECT 195.675 -13.765 196.005 -13.435 ;
        RECT 194.315 -13.765 194.645 -13.435 ;
        RECT 192.955 -13.765 193.285 -13.435 ;
        RECT 191.595 -13.765 191.925 -13.435 ;
        RECT 190.235 -13.765 190.565 -13.435 ;
        RECT 188.875 -13.765 189.205 -13.435 ;
        RECT 187.515 -13.765 187.845 -13.435 ;
        RECT 186.155 -13.765 186.485 -13.435 ;
        RECT 184.795 -13.765 185.125 -13.435 ;
        RECT 183.435 -13.765 183.765 -13.435 ;
        RECT 182.075 -13.765 182.405 -13.435 ;
        RECT 180.715 -13.765 181.045 -13.435 ;
        RECT 179.355 -13.765 179.685 -13.435 ;
        RECT 177.995 -13.765 178.325 -13.435 ;
        RECT 176.635 -13.765 176.965 -13.435 ;
        RECT 175.275 -13.765 175.605 -13.435 ;
        RECT 173.915 -13.765 174.245 -13.435 ;
        RECT 172.555 -13.765 172.885 -13.435 ;
        RECT 171.195 -13.765 171.525 -13.435 ;
        RECT 169.835 -13.765 170.165 -13.435 ;
        RECT 168.475 -13.765 168.805 -13.435 ;
        RECT 167.115 -13.765 167.445 -13.435 ;
        RECT 165.755 -13.765 166.085 -13.435 ;
        RECT 164.395 -13.765 164.725 -13.435 ;
        RECT 163.035 -13.765 163.365 -13.435 ;
        RECT 161.675 -13.765 162.005 -13.435 ;
        RECT 160.315 -13.765 160.645 -13.435 ;
        RECT 158.955 -13.765 159.285 -13.435 ;
        RECT 157.595 -13.765 157.925 -13.435 ;
        RECT 156.235 -13.765 156.565 -13.435 ;
        RECT 154.875 -13.765 155.205 -13.435 ;
        RECT 153.515 -13.765 153.845 -13.435 ;
        RECT 152.155 -13.765 152.485 -13.435 ;
        RECT 150.795 -13.765 151.125 -13.435 ;
        RECT 149.435 -13.765 149.765 -13.435 ;
        RECT 148.075 -13.765 148.405 -13.435 ;
        RECT 146.715 -13.765 147.045 -13.435 ;
        RECT 145.355 -13.765 145.685 -13.435 ;
        RECT 143.995 -13.765 144.325 -13.435 ;
        RECT 142.635 -13.765 142.965 -13.435 ;
        RECT 141.275 -13.765 141.605 -13.435 ;
        RECT 139.915 -13.765 140.245 -13.435 ;
        RECT 138.555 -13.765 138.885 -13.435 ;
        RECT 137.195 -13.765 137.525 -13.435 ;
        RECT 135.835 -13.765 136.165 -13.435 ;
        RECT 134.475 -13.765 134.805 -13.435 ;
        RECT 133.115 -13.765 133.445 -13.435 ;
        RECT 131.755 -13.765 132.085 -13.435 ;
        RECT 130.395 -13.765 130.725 -13.435 ;
        RECT 129.035 -13.765 129.365 -13.435 ;
        RECT 127.675 -13.765 128.005 -13.435 ;
        RECT 126.315 -13.765 126.645 -13.435 ;
        RECT 124.955 -13.765 125.285 -13.435 ;
        RECT 123.595 -13.765 123.925 -13.435 ;
        RECT 122.235 -13.765 122.565 -13.435 ;
        RECT 120.875 -13.765 121.205 -13.435 ;
        RECT 119.515 -13.765 119.845 -13.435 ;
        RECT 118.155 -13.765 118.485 -13.435 ;
        RECT 116.795 -13.765 117.125 -13.435 ;
        RECT 115.435 -13.765 115.765 -13.435 ;
        RECT 114.075 -13.765 114.405 -13.435 ;
        RECT 112.715 -13.765 113.045 -13.435 ;
        RECT 111.355 -13.765 111.685 -13.435 ;
        RECT 109.995 -13.765 110.325 -13.435 ;
        RECT 108.635 -13.765 108.965 -13.435 ;
        RECT 107.275 -13.765 107.605 -13.435 ;
        RECT 105.915 -13.765 106.245 -13.435 ;
        RECT 104.555 -13.765 104.885 -13.435 ;
        RECT 103.195 -13.765 103.525 -13.435 ;
        RECT 101.835 -13.765 102.165 -13.435 ;
        RECT 100.475 -13.765 100.805 -13.435 ;
        RECT 99.115 -13.765 99.445 -13.435 ;
        RECT 97.755 -13.765 98.085 -13.435 ;
        RECT 96.395 -13.765 96.725 -13.435 ;
        RECT 95.035 -13.765 95.365 -13.435 ;
        RECT 93.675 -13.765 94.005 -13.435 ;
        RECT 92.315 -13.765 92.645 -13.435 ;
        RECT 90.955 -13.765 91.285 -13.435 ;
        RECT 89.595 -13.765 89.925 -13.435 ;
        RECT 88.235 -13.765 88.565 -13.435 ;
        RECT 86.875 -13.765 87.205 -13.435 ;
        RECT 85.515 -13.765 85.845 -13.435 ;
        RECT 84.155 -13.765 84.485 -13.435 ;
        RECT 82.795 -13.765 83.125 -13.435 ;
        RECT 81.435 -13.765 81.765 -13.435 ;
        RECT 80.075 -13.765 80.405 -13.435 ;
        RECT 78.715 -13.765 79.045 -13.435 ;
        RECT 77.355 -13.765 77.685 -13.435 ;
        RECT 75.995 -13.765 76.325 -13.435 ;
        RECT 74.635 -13.765 74.965 -13.435 ;
        RECT 73.275 -13.765 73.605 -13.435 ;
        RECT 71.915 -13.765 72.245 -13.435 ;
        RECT 70.555 -13.765 70.885 -13.435 ;
        RECT 69.195 -13.765 69.525 -13.435 ;
        RECT 67.835 -13.765 68.165 -13.435 ;
        RECT 66.475 -13.765 66.805 -13.435 ;
        RECT 65.115 -13.765 65.445 -13.435 ;
        RECT 63.755 -13.765 64.085 -13.435 ;
        RECT 62.395 -13.765 62.725 -13.435 ;
        RECT 61.035 -13.765 61.365 -13.435 ;
        RECT 59.675 -13.765 60.005 -13.435 ;
        RECT 58.315 -13.765 58.645 -13.435 ;
        RECT 56.955 -13.765 57.285 -13.435 ;
        RECT 55.595 -13.765 55.925 -13.435 ;
        RECT 54.235 -13.765 54.565 -13.435 ;
        RECT 52.875 -13.765 53.205 -13.435 ;
        RECT 51.515 -13.765 51.845 -13.435 ;
        RECT 50.155 -13.765 50.485 -13.435 ;
        RECT 48.795 -13.765 49.125 -13.435 ;
        RECT 47.435 -13.765 47.765 -13.435 ;
        RECT 46.075 -13.765 46.405 -13.435 ;
        RECT 44.715 -13.765 45.045 -13.435 ;
        RECT 43.355 -13.765 43.685 -13.435 ;
        RECT 41.995 -13.765 42.325 -13.435 ;
        RECT 40.635 -13.765 40.965 -13.435 ;
        RECT 39.275 -13.765 39.605 -13.435 ;
        RECT 37.915 -13.765 38.245 -13.435 ;
        RECT 36.555 -13.765 36.885 -13.435 ;
        RECT 35.195 -13.765 35.525 -13.435 ;
        RECT 33.835 -13.765 34.165 -13.435 ;
        RECT 32.475 -13.765 32.805 -13.435 ;
        RECT 31.115 -13.765 31.445 -13.435 ;
        RECT 29.755 -13.765 30.085 -13.435 ;
        RECT 28.395 -13.765 28.725 -13.435 ;
        RECT 27.035 -13.765 27.365 -13.435 ;
        RECT 25.675 -13.765 26.005 -13.435 ;
        RECT 24.315 -13.765 24.645 -13.435 ;
        RECT 22.955 -13.765 23.285 -13.435 ;
        RECT 21.595 -13.765 21.925 -13.435 ;
        RECT 20.235 -13.765 20.565 -13.435 ;
        RECT 18.875 -13.765 19.205 -13.435 ;
        RECT 17.515 -13.765 17.845 -13.435 ;
        RECT 16.155 -13.765 16.485 -13.435 ;
        RECT 14.795 -13.765 15.125 -13.435 ;
        RECT 13.435 -13.765 13.765 -13.435 ;
        RECT 12.075 -13.765 12.405 -13.435 ;
        RECT 10.715 -13.765 11.045 -13.435 ;
        RECT 9.355 -13.765 9.685 -13.435 ;
        RECT 7.995 -13.765 8.325 -13.435 ;
        RECT 6.635 -13.765 6.965 -13.435 ;
        RECT 5.275 -13.765 5.605 -13.435 ;
        RECT 3.915 -13.765 4.245 -13.435 ;
        RECT 2.555 -13.765 2.885 -13.435 ;
        RECT 1.195 -13.765 1.525 -13.435 ;
        RECT -0.165 -13.765 0.165 -13.435 ;
        RECT -1.525 -13.765 -1.195 -13.435 ;
        RECT -1.525 -13.76 678.475 -13.44 ;
        RECT 677.115 -13.765 677.445 -13.435 ;
        RECT 675.755 -13.765 676.085 -13.435 ;
        RECT 674.395 -13.765 674.725 -13.435 ;
        RECT 673.035 -13.765 673.365 -13.435 ;
        RECT 671.675 -13.765 672.005 -13.435 ;
        RECT 670.315 -13.765 670.645 -13.435 ;
        RECT 668.955 -13.765 669.285 -13.435 ;
        RECT 667.595 -13.765 667.925 -13.435 ;
        RECT 666.235 -13.765 666.565 -13.435 ;
        RECT 664.875 -13.765 665.205 -13.435 ;
        RECT 663.515 -13.765 663.845 -13.435 ;
        RECT 662.155 -13.765 662.485 -13.435 ;
        RECT 660.795 -13.765 661.125 -13.435 ;
        RECT 659.435 -13.765 659.765 -13.435 ;
        RECT 658.075 -13.765 658.405 -13.435 ;
        RECT 656.715 -13.765 657.045 -13.435 ;
        RECT 655.355 -13.765 655.685 -13.435 ;
        RECT 653.995 -13.765 654.325 -13.435 ;
        RECT 652.635 -13.765 652.965 -13.435 ;
        RECT 651.275 -13.765 651.605 -13.435 ;
        RECT 649.915 -13.765 650.245 -13.435 ;
        RECT 648.555 -13.765 648.885 -13.435 ;
        RECT 647.195 -13.765 647.525 -13.435 ;
        RECT 954.555 -13.765 954.885 -13.435 ;
        RECT 678.475 -13.76 954.885 -13.44 ;
        RECT 953.195 -13.765 953.525 -13.435 ;
        RECT 951.835 -13.765 952.165 -13.435 ;
        RECT 950.475 -13.765 950.805 -13.435 ;
        RECT 949.115 -13.765 949.445 -13.435 ;
        RECT 947.755 -13.765 948.085 -13.435 ;
        RECT 946.395 -13.765 946.725 -13.435 ;
        RECT 945.035 -13.765 945.365 -13.435 ;
        RECT 943.675 -13.765 944.005 -13.435 ;
        RECT 942.315 -13.765 942.645 -13.435 ;
        RECT 940.955 -13.765 941.285 -13.435 ;
        RECT 939.595 -13.765 939.925 -13.435 ;
        RECT 938.235 -13.765 938.565 -13.435 ;
        RECT 936.875 -13.765 937.205 -13.435 ;
        RECT 935.515 -13.765 935.845 -13.435 ;
        RECT 934.155 -13.765 934.485 -13.435 ;
        RECT 932.795 -13.765 933.125 -13.435 ;
        RECT 931.435 -13.765 931.765 -13.435 ;
        RECT 930.075 -13.765 930.405 -13.435 ;
        RECT 928.715 -13.765 929.045 -13.435 ;
        RECT 927.355 -13.765 927.685 -13.435 ;
        RECT 925.995 -13.765 926.325 -13.435 ;
        RECT 924.635 -13.765 924.965 -13.435 ;
        RECT 923.275 -13.765 923.605 -13.435 ;
        RECT 921.915 -13.765 922.245 -13.435 ;
        RECT 920.555 -13.765 920.885 -13.435 ;
        RECT 919.195 -13.765 919.525 -13.435 ;
        RECT 917.835 -13.765 918.165 -13.435 ;
        RECT 916.475 -13.765 916.805 -13.435 ;
        RECT 915.115 -13.765 915.445 -13.435 ;
        RECT 913.755 -13.765 914.085 -13.435 ;
        RECT 912.395 -13.765 912.725 -13.435 ;
        RECT 911.035 -13.765 911.365 -13.435 ;
        RECT 909.675 -13.765 910.005 -13.435 ;
        RECT 908.315 -13.765 908.645 -13.435 ;
        RECT 906.955 -13.765 907.285 -13.435 ;
        RECT 905.595 -13.765 905.925 -13.435 ;
        RECT 904.235 -13.765 904.565 -13.435 ;
        RECT 902.875 -13.765 903.205 -13.435 ;
        RECT 901.515 -13.765 901.845 -13.435 ;
        RECT 900.155 -13.765 900.485 -13.435 ;
        RECT 898.795 -13.765 899.125 -13.435 ;
        RECT 897.435 -13.765 897.765 -13.435 ;
        RECT 896.075 -13.765 896.405 -13.435 ;
        RECT 894.715 -13.765 895.045 -13.435 ;
        RECT 893.355 -13.765 893.685 -13.435 ;
        RECT 891.995 -13.765 892.325 -13.435 ;
        RECT 890.635 -13.765 890.965 -13.435 ;
        RECT 889.275 -13.765 889.605 -13.435 ;
        RECT 887.915 -13.765 888.245 -13.435 ;
        RECT 886.555 -13.765 886.885 -13.435 ;
        RECT 885.195 -13.765 885.525 -13.435 ;
        RECT 883.835 -13.765 884.165 -13.435 ;
        RECT 882.475 -13.765 882.805 -13.435 ;
        RECT 881.115 -13.765 881.445 -13.435 ;
        RECT 879.755 -13.765 880.085 -13.435 ;
        RECT 878.395 -13.765 878.725 -13.435 ;
        RECT 877.035 -13.765 877.365 -13.435 ;
        RECT 875.675 -13.765 876.005 -13.435 ;
        RECT 874.315 -13.765 874.645 -13.435 ;
        RECT 872.955 -13.765 873.285 -13.435 ;
        RECT 871.595 -13.765 871.925 -13.435 ;
        RECT 870.235 -13.765 870.565 -13.435 ;
        RECT 868.875 -13.765 869.205 -13.435 ;
        RECT 867.515 -13.765 867.845 -13.435 ;
        RECT 866.155 -13.765 866.485 -13.435 ;
        RECT 864.795 -13.765 865.125 -13.435 ;
        RECT 863.435 -13.765 863.765 -13.435 ;
        RECT 862.075 -13.765 862.405 -13.435 ;
        RECT 860.715 -13.765 861.045 -13.435 ;
        RECT 859.355 -13.765 859.685 -13.435 ;
        RECT 857.995 -13.765 858.325 -13.435 ;
        RECT 856.635 -13.765 856.965 -13.435 ;
        RECT 855.275 -13.765 855.605 -13.435 ;
        RECT 853.915 -13.765 854.245 -13.435 ;
        RECT 852.555 -13.765 852.885 -13.435 ;
        RECT 851.195 -13.765 851.525 -13.435 ;
        RECT 849.835 -13.765 850.165 -13.435 ;
        RECT 848.475 -13.765 848.805 -13.435 ;
        RECT 847.115 -13.765 847.445 -13.435 ;
        RECT 845.755 -13.765 846.085 -13.435 ;
        RECT 844.395 -13.765 844.725 -13.435 ;
        RECT 843.035 -13.765 843.365 -13.435 ;
        RECT 841.675 -13.765 842.005 -13.435 ;
        RECT 840.315 -13.765 840.645 -13.435 ;
        RECT 838.955 -13.765 839.285 -13.435 ;
        RECT 837.595 -13.765 837.925 -13.435 ;
        RECT 836.235 -13.765 836.565 -13.435 ;
        RECT 834.875 -13.765 835.205 -13.435 ;
        RECT 833.515 -13.765 833.845 -13.435 ;
        RECT 832.155 -13.765 832.485 -13.435 ;
        RECT 830.795 -13.765 831.125 -13.435 ;
        RECT 829.435 -13.765 829.765 -13.435 ;
        RECT 828.075 -13.765 828.405 -13.435 ;
        RECT 826.715 -13.765 827.045 -13.435 ;
        RECT 825.355 -13.765 825.685 -13.435 ;
        RECT 823.995 -13.765 824.325 -13.435 ;
        RECT 822.635 -13.765 822.965 -13.435 ;
        RECT 821.275 -13.765 821.605 -13.435 ;
        RECT 819.915 -13.765 820.245 -13.435 ;
        RECT 818.555 -13.765 818.885 -13.435 ;
        RECT 817.195 -13.765 817.525 -13.435 ;
        RECT 815.835 -13.765 816.165 -13.435 ;
        RECT 814.475 -13.765 814.805 -13.435 ;
        RECT 813.115 -13.765 813.445 -13.435 ;
        RECT 811.755 -13.765 812.085 -13.435 ;
        RECT 810.395 -13.765 810.725 -13.435 ;
        RECT 809.035 -13.765 809.365 -13.435 ;
        RECT 807.675 -13.765 808.005 -13.435 ;
        RECT 806.315 -13.765 806.645 -13.435 ;
        RECT 804.955 -13.765 805.285 -13.435 ;
        RECT 803.595 -13.765 803.925 -13.435 ;
        RECT 802.235 -13.765 802.565 -13.435 ;
        RECT 800.875 -13.765 801.205 -13.435 ;
        RECT 799.515 -13.765 799.845 -13.435 ;
        RECT 798.155 -13.765 798.485 -13.435 ;
        RECT 796.795 -13.765 797.125 -13.435 ;
        RECT 795.435 -13.765 795.765 -13.435 ;
        RECT 794.075 -13.765 794.405 -13.435 ;
        RECT 792.715 -13.765 793.045 -13.435 ;
        RECT 791.355 -13.765 791.685 -13.435 ;
        RECT 789.995 -13.765 790.325 -13.435 ;
        RECT 788.635 -13.765 788.965 -13.435 ;
        RECT 787.275 -13.765 787.605 -13.435 ;
        RECT 785.915 -13.765 786.245 -13.435 ;
        RECT 784.555 -13.765 784.885 -13.435 ;
        RECT 783.195 -13.765 783.525 -13.435 ;
        RECT 781.835 -13.765 782.165 -13.435 ;
        RECT 780.475 -13.765 780.805 -13.435 ;
        RECT 779.115 -13.765 779.445 -13.435 ;
        RECT 777.755 -13.765 778.085 -13.435 ;
        RECT 776.395 -13.765 776.725 -13.435 ;
        RECT 775.035 -13.765 775.365 -13.435 ;
        RECT 773.675 -13.765 774.005 -13.435 ;
        RECT 772.315 -13.765 772.645 -13.435 ;
        RECT 770.955 -13.765 771.285 -13.435 ;
        RECT 769.595 -13.765 769.925 -13.435 ;
        RECT 768.235 -13.765 768.565 -13.435 ;
        RECT 766.875 -13.765 767.205 -13.435 ;
        RECT 765.515 -13.765 765.845 -13.435 ;
        RECT 764.155 -13.765 764.485 -13.435 ;
        RECT 762.795 -13.765 763.125 -13.435 ;
        RECT 761.435 -13.765 761.765 -13.435 ;
        RECT 760.075 -13.765 760.405 -13.435 ;
        RECT 758.715 -13.765 759.045 -13.435 ;
        RECT 757.355 -13.765 757.685 -13.435 ;
        RECT 755.995 -13.765 756.325 -13.435 ;
        RECT 754.635 -13.765 754.965 -13.435 ;
        RECT 753.275 -13.765 753.605 -13.435 ;
        RECT 751.915 -13.765 752.245 -13.435 ;
        RECT 750.555 -13.765 750.885 -13.435 ;
        RECT 749.195 -13.765 749.525 -13.435 ;
        RECT 747.835 -13.765 748.165 -13.435 ;
        RECT 746.475 -13.765 746.805 -13.435 ;
        RECT 745.115 -13.765 745.445 -13.435 ;
        RECT 743.755 -13.765 744.085 -13.435 ;
        RECT 742.395 -13.765 742.725 -13.435 ;
        RECT 741.035 -13.765 741.365 -13.435 ;
        RECT 739.675 -13.765 740.005 -13.435 ;
        RECT 738.315 -13.765 738.645 -13.435 ;
        RECT 736.955 -13.765 737.285 -13.435 ;
        RECT 735.595 -13.765 735.925 -13.435 ;
        RECT 734.235 -13.765 734.565 -13.435 ;
        RECT 732.875 -13.765 733.205 -13.435 ;
        RECT 731.515 -13.765 731.845 -13.435 ;
        RECT 730.155 -13.765 730.485 -13.435 ;
        RECT 728.795 -13.765 729.125 -13.435 ;
        RECT 727.435 -13.765 727.765 -13.435 ;
        RECT 726.075 -13.765 726.405 -13.435 ;
        RECT 724.715 -13.765 725.045 -13.435 ;
        RECT 723.355 -13.765 723.685 -13.435 ;
        RECT 721.995 -13.765 722.325 -13.435 ;
        RECT 720.635 -13.765 720.965 -13.435 ;
        RECT 719.275 -13.765 719.605 -13.435 ;
        RECT 717.915 -13.765 718.245 -13.435 ;
        RECT 716.555 -13.765 716.885 -13.435 ;
        RECT 715.195 -13.765 715.525 -13.435 ;
        RECT 713.835 -13.765 714.165 -13.435 ;
        RECT 712.475 -13.765 712.805 -13.435 ;
        RECT 711.115 -13.765 711.445 -13.435 ;
        RECT 709.755 -13.765 710.085 -13.435 ;
        RECT 708.395 -13.765 708.725 -13.435 ;
        RECT 707.035 -13.765 707.365 -13.435 ;
        RECT 705.675 -13.765 706.005 -13.435 ;
        RECT 704.315 -13.765 704.645 -13.435 ;
        RECT 702.955 -13.765 703.285 -13.435 ;
        RECT 701.595 -13.765 701.925 -13.435 ;
        RECT 700.235 -13.765 700.565 -13.435 ;
        RECT 698.875 -13.765 699.205 -13.435 ;
        RECT 697.515 -13.765 697.845 -13.435 ;
        RECT 696.155 -13.765 696.485 -13.435 ;
        RECT 694.795 -13.765 695.125 -13.435 ;
        RECT 693.435 -13.765 693.765 -13.435 ;
        RECT 692.075 -13.765 692.405 -13.435 ;
        RECT 690.715 -13.765 691.045 -13.435 ;
        RECT 689.355 -13.765 689.685 -13.435 ;
        RECT 687.995 -13.765 688.325 -13.435 ;
        RECT 686.635 -13.765 686.965 -13.435 ;
        RECT 685.275 -13.765 685.605 -13.435 ;
        RECT 683.915 -13.765 684.245 -13.435 ;
        RECT 682.555 -13.765 682.885 -13.435 ;
        RECT 681.195 -13.765 681.525 -13.435 ;
        RECT 679.835 -13.765 680.165 -13.435 ;
        RECT 678.475 -13.765 678.805 -13.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -9.68 678.475 -9.36 ;
        RECT 677.115 -9.685 677.445 -9.355 ;
        RECT 675.755 -9.685 676.085 -9.355 ;
        RECT 674.395 -9.685 674.725 -9.355 ;
        RECT 673.035 -9.685 673.365 -9.355 ;
        RECT 671.675 -9.685 672.005 -9.355 ;
        RECT 670.315 -9.685 670.645 -9.355 ;
        RECT 668.955 -9.685 669.285 -9.355 ;
        RECT 667.595 -9.685 667.925 -9.355 ;
        RECT 666.235 -9.685 666.565 -9.355 ;
        RECT 664.875 -9.685 665.205 -9.355 ;
        RECT 663.515 -9.685 663.845 -9.355 ;
        RECT 662.155 -9.685 662.485 -9.355 ;
        RECT 660.795 -9.685 661.125 -9.355 ;
        RECT 659.435 -9.685 659.765 -9.355 ;
        RECT 658.075 -9.685 658.405 -9.355 ;
        RECT 656.715 -9.685 657.045 -9.355 ;
        RECT 655.355 -9.685 655.685 -9.355 ;
        RECT 653.995 -9.685 654.325 -9.355 ;
        RECT 652.635 -9.685 652.965 -9.355 ;
        RECT 651.275 -9.685 651.605 -9.355 ;
        RECT 649.915 -9.685 650.245 -9.355 ;
        RECT 648.555 -9.685 648.885 -9.355 ;
        RECT 647.195 -9.685 647.525 -9.355 ;
        RECT 645.835 -9.685 646.165 -9.355 ;
        RECT 644.475 -9.685 644.805 -9.355 ;
        RECT 643.115 -9.685 643.445 -9.355 ;
        RECT 641.755 -9.685 642.085 -9.355 ;
        RECT 640.395 -9.685 640.725 -9.355 ;
        RECT 639.035 -9.685 639.365 -9.355 ;
        RECT 637.675 -9.685 638.005 -9.355 ;
        RECT 636.315 -9.685 636.645 -9.355 ;
        RECT 634.955 -9.685 635.285 -9.355 ;
        RECT 633.595 -9.685 633.925 -9.355 ;
        RECT 632.235 -9.685 632.565 -9.355 ;
        RECT 630.875 -9.685 631.205 -9.355 ;
        RECT 629.515 -9.685 629.845 -9.355 ;
        RECT 628.155 -9.685 628.485 -9.355 ;
        RECT 626.795 -9.685 627.125 -9.355 ;
        RECT 625.435 -9.685 625.765 -9.355 ;
        RECT 624.075 -9.685 624.405 -9.355 ;
        RECT 622.715 -9.685 623.045 -9.355 ;
        RECT 621.355 -9.685 621.685 -9.355 ;
        RECT 619.995 -9.685 620.325 -9.355 ;
        RECT 618.635 -9.685 618.965 -9.355 ;
        RECT 617.275 -9.685 617.605 -9.355 ;
        RECT 615.915 -9.685 616.245 -9.355 ;
        RECT 614.555 -9.685 614.885 -9.355 ;
        RECT 613.195 -9.685 613.525 -9.355 ;
        RECT 611.835 -9.685 612.165 -9.355 ;
        RECT 610.475 -9.685 610.805 -9.355 ;
        RECT 609.115 -9.685 609.445 -9.355 ;
        RECT 607.755 -9.685 608.085 -9.355 ;
        RECT 606.395 -9.685 606.725 -9.355 ;
        RECT 605.035 -9.685 605.365 -9.355 ;
        RECT 603.675 -9.685 604.005 -9.355 ;
        RECT 602.315 -9.685 602.645 -9.355 ;
        RECT 600.955 -9.685 601.285 -9.355 ;
        RECT 599.595 -9.685 599.925 -9.355 ;
        RECT 598.235 -9.685 598.565 -9.355 ;
        RECT 596.875 -9.685 597.205 -9.355 ;
        RECT 595.515 -9.685 595.845 -9.355 ;
        RECT 594.155 -9.685 594.485 -9.355 ;
        RECT 592.795 -9.685 593.125 -9.355 ;
        RECT 591.435 -9.685 591.765 -9.355 ;
        RECT 590.075 -9.685 590.405 -9.355 ;
        RECT 588.715 -9.685 589.045 -9.355 ;
        RECT 587.355 -9.685 587.685 -9.355 ;
        RECT 585.995 -9.685 586.325 -9.355 ;
        RECT 584.635 -9.685 584.965 -9.355 ;
        RECT 583.275 -9.685 583.605 -9.355 ;
        RECT 581.915 -9.685 582.245 -9.355 ;
        RECT 580.555 -9.685 580.885 -9.355 ;
        RECT 579.195 -9.685 579.525 -9.355 ;
        RECT 577.835 -9.685 578.165 -9.355 ;
        RECT 576.475 -9.685 576.805 -9.355 ;
        RECT 575.115 -9.685 575.445 -9.355 ;
        RECT 573.755 -9.685 574.085 -9.355 ;
        RECT 572.395 -9.685 572.725 -9.355 ;
        RECT 571.035 -9.685 571.365 -9.355 ;
        RECT 569.675 -9.685 570.005 -9.355 ;
        RECT 568.315 -9.685 568.645 -9.355 ;
        RECT 566.955 -9.685 567.285 -9.355 ;
        RECT 565.595 -9.685 565.925 -9.355 ;
        RECT 564.235 -9.685 564.565 -9.355 ;
        RECT 562.875 -9.685 563.205 -9.355 ;
        RECT 561.515 -9.685 561.845 -9.355 ;
        RECT 560.155 -9.685 560.485 -9.355 ;
        RECT 558.795 -9.685 559.125 -9.355 ;
        RECT 557.435 -9.685 557.765 -9.355 ;
        RECT 556.075 -9.685 556.405 -9.355 ;
        RECT 554.715 -9.685 555.045 -9.355 ;
        RECT 553.355 -9.685 553.685 -9.355 ;
        RECT 551.995 -9.685 552.325 -9.355 ;
        RECT 550.635 -9.685 550.965 -9.355 ;
        RECT 549.275 -9.685 549.605 -9.355 ;
        RECT 547.915 -9.685 548.245 -9.355 ;
        RECT 546.555 -9.685 546.885 -9.355 ;
        RECT 545.195 -9.685 545.525 -9.355 ;
        RECT 543.835 -9.685 544.165 -9.355 ;
        RECT 542.475 -9.685 542.805 -9.355 ;
        RECT 541.115 -9.685 541.445 -9.355 ;
        RECT 539.755 -9.685 540.085 -9.355 ;
        RECT 538.395 -9.685 538.725 -9.355 ;
        RECT 537.035 -9.685 537.365 -9.355 ;
        RECT 535.675 -9.685 536.005 -9.355 ;
        RECT 534.315 -9.685 534.645 -9.355 ;
        RECT 532.955 -9.685 533.285 -9.355 ;
        RECT 531.595 -9.685 531.925 -9.355 ;
        RECT 530.235 -9.685 530.565 -9.355 ;
        RECT 528.875 -9.685 529.205 -9.355 ;
        RECT 527.515 -9.685 527.845 -9.355 ;
        RECT 526.155 -9.685 526.485 -9.355 ;
        RECT 524.795 -9.685 525.125 -9.355 ;
        RECT 523.435 -9.685 523.765 -9.355 ;
        RECT 522.075 -9.685 522.405 -9.355 ;
        RECT 520.715 -9.685 521.045 -9.355 ;
        RECT 519.355 -9.685 519.685 -9.355 ;
        RECT 517.995 -9.685 518.325 -9.355 ;
        RECT 516.635 -9.685 516.965 -9.355 ;
        RECT 515.275 -9.685 515.605 -9.355 ;
        RECT 513.915 -9.685 514.245 -9.355 ;
        RECT 512.555 -9.685 512.885 -9.355 ;
        RECT 511.195 -9.685 511.525 -9.355 ;
        RECT 509.835 -9.685 510.165 -9.355 ;
        RECT 508.475 -9.685 508.805 -9.355 ;
        RECT 507.115 -9.685 507.445 -9.355 ;
        RECT 505.755 -9.685 506.085 -9.355 ;
        RECT 504.395 -9.685 504.725 -9.355 ;
        RECT 503.035 -9.685 503.365 -9.355 ;
        RECT 501.675 -9.685 502.005 -9.355 ;
        RECT 500.315 -9.685 500.645 -9.355 ;
        RECT 498.955 -9.685 499.285 -9.355 ;
        RECT 497.595 -9.685 497.925 -9.355 ;
        RECT 496.235 -9.685 496.565 -9.355 ;
        RECT 494.875 -9.685 495.205 -9.355 ;
        RECT 493.515 -9.685 493.845 -9.355 ;
        RECT 492.155 -9.685 492.485 -9.355 ;
        RECT 490.795 -9.685 491.125 -9.355 ;
        RECT 489.435 -9.685 489.765 -9.355 ;
        RECT 488.075 -9.685 488.405 -9.355 ;
        RECT 486.715 -9.685 487.045 -9.355 ;
        RECT 485.355 -9.685 485.685 -9.355 ;
        RECT 483.995 -9.685 484.325 -9.355 ;
        RECT 482.635 -9.685 482.965 -9.355 ;
        RECT 481.275 -9.685 481.605 -9.355 ;
        RECT 479.915 -9.685 480.245 -9.355 ;
        RECT 478.555 -9.685 478.885 -9.355 ;
        RECT 477.195 -9.685 477.525 -9.355 ;
        RECT 475.835 -9.685 476.165 -9.355 ;
        RECT 474.475 -9.685 474.805 -9.355 ;
        RECT 473.115 -9.685 473.445 -9.355 ;
        RECT 471.755 -9.685 472.085 -9.355 ;
        RECT 470.395 -9.685 470.725 -9.355 ;
        RECT 469.035 -9.685 469.365 -9.355 ;
        RECT 467.675 -9.685 468.005 -9.355 ;
        RECT 466.315 -9.685 466.645 -9.355 ;
        RECT 464.955 -9.685 465.285 -9.355 ;
        RECT 463.595 -9.685 463.925 -9.355 ;
        RECT 462.235 -9.685 462.565 -9.355 ;
        RECT 460.875 -9.685 461.205 -9.355 ;
        RECT 459.515 -9.685 459.845 -9.355 ;
        RECT 458.155 -9.685 458.485 -9.355 ;
        RECT 456.795 -9.685 457.125 -9.355 ;
        RECT 455.435 -9.685 455.765 -9.355 ;
        RECT 454.075 -9.685 454.405 -9.355 ;
        RECT 452.715 -9.685 453.045 -9.355 ;
        RECT 451.355 -9.685 451.685 -9.355 ;
        RECT 449.995 -9.685 450.325 -9.355 ;
        RECT 448.635 -9.685 448.965 -9.355 ;
        RECT 447.275 -9.685 447.605 -9.355 ;
        RECT 445.915 -9.685 446.245 -9.355 ;
        RECT 444.555 -9.685 444.885 -9.355 ;
        RECT 443.195 -9.685 443.525 -9.355 ;
        RECT 441.835 -9.685 442.165 -9.355 ;
        RECT 440.475 -9.685 440.805 -9.355 ;
        RECT 439.115 -9.685 439.445 -9.355 ;
        RECT 437.755 -9.685 438.085 -9.355 ;
        RECT 436.395 -9.685 436.725 -9.355 ;
        RECT 435.035 -9.685 435.365 -9.355 ;
        RECT 433.675 -9.685 434.005 -9.355 ;
        RECT 432.315 -9.685 432.645 -9.355 ;
        RECT 430.955 -9.685 431.285 -9.355 ;
        RECT 429.595 -9.685 429.925 -9.355 ;
        RECT 428.235 -9.685 428.565 -9.355 ;
        RECT 426.875 -9.685 427.205 -9.355 ;
        RECT 425.515 -9.685 425.845 -9.355 ;
        RECT 424.155 -9.685 424.485 -9.355 ;
        RECT 422.795 -9.685 423.125 -9.355 ;
        RECT 421.435 -9.685 421.765 -9.355 ;
        RECT 420.075 -9.685 420.405 -9.355 ;
        RECT 418.715 -9.685 419.045 -9.355 ;
        RECT 417.355 -9.685 417.685 -9.355 ;
        RECT 415.995 -9.685 416.325 -9.355 ;
        RECT 414.635 -9.685 414.965 -9.355 ;
        RECT 413.275 -9.685 413.605 -9.355 ;
        RECT 411.915 -9.685 412.245 -9.355 ;
        RECT 410.555 -9.685 410.885 -9.355 ;
        RECT 409.195 -9.685 409.525 -9.355 ;
        RECT 407.835 -9.685 408.165 -9.355 ;
        RECT 406.475 -9.685 406.805 -9.355 ;
        RECT 405.115 -9.685 405.445 -9.355 ;
        RECT 403.755 -9.685 404.085 -9.355 ;
        RECT 402.395 -9.685 402.725 -9.355 ;
        RECT 401.035 -9.685 401.365 -9.355 ;
        RECT 399.675 -9.685 400.005 -9.355 ;
        RECT 398.315 -9.685 398.645 -9.355 ;
        RECT 396.955 -9.685 397.285 -9.355 ;
        RECT 395.595 -9.685 395.925 -9.355 ;
        RECT 394.235 -9.685 394.565 -9.355 ;
        RECT 392.875 -9.685 393.205 -9.355 ;
        RECT 391.515 -9.685 391.845 -9.355 ;
        RECT 390.155 -9.685 390.485 -9.355 ;
        RECT 388.795 -9.685 389.125 -9.355 ;
        RECT 387.435 -9.685 387.765 -9.355 ;
        RECT 386.075 -9.685 386.405 -9.355 ;
        RECT 384.715 -9.685 385.045 -9.355 ;
        RECT 383.355 -9.685 383.685 -9.355 ;
        RECT 381.995 -9.685 382.325 -9.355 ;
        RECT 380.635 -9.685 380.965 -9.355 ;
        RECT 379.275 -9.685 379.605 -9.355 ;
        RECT 377.915 -9.685 378.245 -9.355 ;
        RECT 376.555 -9.685 376.885 -9.355 ;
        RECT 375.195 -9.685 375.525 -9.355 ;
        RECT 373.835 -9.685 374.165 -9.355 ;
        RECT 372.475 -9.685 372.805 -9.355 ;
        RECT 371.115 -9.685 371.445 -9.355 ;
        RECT 369.755 -9.685 370.085 -9.355 ;
        RECT 368.395 -9.685 368.725 -9.355 ;
        RECT 367.035 -9.685 367.365 -9.355 ;
        RECT 365.675 -9.685 366.005 -9.355 ;
        RECT 364.315 -9.685 364.645 -9.355 ;
        RECT 362.955 -9.685 363.285 -9.355 ;
        RECT 361.595 -9.685 361.925 -9.355 ;
        RECT 360.235 -9.685 360.565 -9.355 ;
        RECT 358.875 -9.685 359.205 -9.355 ;
        RECT 357.515 -9.685 357.845 -9.355 ;
        RECT 356.155 -9.685 356.485 -9.355 ;
        RECT 354.795 -9.685 355.125 -9.355 ;
        RECT 353.435 -9.685 353.765 -9.355 ;
        RECT 352.075 -9.685 352.405 -9.355 ;
        RECT 350.715 -9.685 351.045 -9.355 ;
        RECT 349.355 -9.685 349.685 -9.355 ;
        RECT 347.995 -9.685 348.325 -9.355 ;
        RECT 346.635 -9.685 346.965 -9.355 ;
        RECT 345.275 -9.685 345.605 -9.355 ;
        RECT 343.915 -9.685 344.245 -9.355 ;
        RECT 342.555 -9.685 342.885 -9.355 ;
        RECT 341.195 -9.685 341.525 -9.355 ;
        RECT 339.835 -9.685 340.165 -9.355 ;
        RECT 338.475 -9.685 338.805 -9.355 ;
        RECT 337.115 -9.685 337.445 -9.355 ;
        RECT 335.755 -9.685 336.085 -9.355 ;
        RECT 334.395 -9.685 334.725 -9.355 ;
        RECT 333.035 -9.685 333.365 -9.355 ;
        RECT 331.675 -9.685 332.005 -9.355 ;
        RECT 330.315 -9.685 330.645 -9.355 ;
        RECT 328.955 -9.685 329.285 -9.355 ;
        RECT 327.595 -9.685 327.925 -9.355 ;
        RECT 326.235 -9.685 326.565 -9.355 ;
        RECT 324.875 -9.685 325.205 -9.355 ;
        RECT 323.515 -9.685 323.845 -9.355 ;
        RECT 322.155 -9.685 322.485 -9.355 ;
        RECT 320.795 -9.685 321.125 -9.355 ;
        RECT 319.435 -9.685 319.765 -9.355 ;
        RECT 318.075 -9.685 318.405 -9.355 ;
        RECT 316.715 -9.685 317.045 -9.355 ;
        RECT 315.355 -9.685 315.685 -9.355 ;
        RECT 313.995 -9.685 314.325 -9.355 ;
        RECT 312.635 -9.685 312.965 -9.355 ;
        RECT 311.275 -9.685 311.605 -9.355 ;
        RECT 309.915 -9.685 310.245 -9.355 ;
        RECT 308.555 -9.685 308.885 -9.355 ;
        RECT 307.195 -9.685 307.525 -9.355 ;
        RECT 305.835 -9.685 306.165 -9.355 ;
        RECT 304.475 -9.685 304.805 -9.355 ;
        RECT 303.115 -9.685 303.445 -9.355 ;
        RECT 301.755 -9.685 302.085 -9.355 ;
        RECT 300.395 -9.685 300.725 -9.355 ;
        RECT 299.035 -9.685 299.365 -9.355 ;
        RECT 297.675 -9.685 298.005 -9.355 ;
        RECT 296.315 -9.685 296.645 -9.355 ;
        RECT 294.955 -9.685 295.285 -9.355 ;
        RECT 293.595 -9.685 293.925 -9.355 ;
        RECT 292.235 -9.685 292.565 -9.355 ;
        RECT 290.875 -9.685 291.205 -9.355 ;
        RECT 289.515 -9.685 289.845 -9.355 ;
        RECT 288.155 -9.685 288.485 -9.355 ;
        RECT 286.795 -9.685 287.125 -9.355 ;
        RECT 285.435 -9.685 285.765 -9.355 ;
        RECT 284.075 -9.685 284.405 -9.355 ;
        RECT 282.715 -9.685 283.045 -9.355 ;
        RECT 281.355 -9.685 281.685 -9.355 ;
        RECT 279.995 -9.685 280.325 -9.355 ;
        RECT 278.635 -9.685 278.965 -9.355 ;
        RECT 277.275 -9.685 277.605 -9.355 ;
        RECT 275.915 -9.685 276.245 -9.355 ;
        RECT 274.555 -9.685 274.885 -9.355 ;
        RECT 273.195 -9.685 273.525 -9.355 ;
        RECT 271.835 -9.685 272.165 -9.355 ;
        RECT 270.475 -9.685 270.805 -9.355 ;
        RECT 269.115 -9.685 269.445 -9.355 ;
        RECT 267.755 -9.685 268.085 -9.355 ;
        RECT 266.395 -9.685 266.725 -9.355 ;
        RECT 265.035 -9.685 265.365 -9.355 ;
        RECT 263.675 -9.685 264.005 -9.355 ;
        RECT 262.315 -9.685 262.645 -9.355 ;
        RECT 260.955 -9.685 261.285 -9.355 ;
        RECT 259.595 -9.685 259.925 -9.355 ;
        RECT 258.235 -9.685 258.565 -9.355 ;
        RECT 256.875 -9.685 257.205 -9.355 ;
        RECT 255.515 -9.685 255.845 -9.355 ;
        RECT 254.155 -9.685 254.485 -9.355 ;
        RECT 252.795 -9.685 253.125 -9.355 ;
        RECT 251.435 -9.685 251.765 -9.355 ;
        RECT 250.075 -9.685 250.405 -9.355 ;
        RECT 248.715 -9.685 249.045 -9.355 ;
        RECT 247.355 -9.685 247.685 -9.355 ;
        RECT 245.995 -9.685 246.325 -9.355 ;
        RECT 244.635 -9.685 244.965 -9.355 ;
        RECT 243.275 -9.685 243.605 -9.355 ;
        RECT 241.915 -9.685 242.245 -9.355 ;
        RECT 240.555 -9.685 240.885 -9.355 ;
        RECT 239.195 -9.685 239.525 -9.355 ;
        RECT 237.835 -9.685 238.165 -9.355 ;
        RECT 236.475 -9.685 236.805 -9.355 ;
        RECT 235.115 -9.685 235.445 -9.355 ;
        RECT 233.755 -9.685 234.085 -9.355 ;
        RECT 232.395 -9.685 232.725 -9.355 ;
        RECT 231.035 -9.685 231.365 -9.355 ;
        RECT 229.675 -9.685 230.005 -9.355 ;
        RECT 228.315 -9.685 228.645 -9.355 ;
        RECT 226.955 -9.685 227.285 -9.355 ;
        RECT 225.595 -9.685 225.925 -9.355 ;
        RECT 224.235 -9.685 224.565 -9.355 ;
        RECT 222.875 -9.685 223.205 -9.355 ;
        RECT 221.515 -9.685 221.845 -9.355 ;
        RECT 220.155 -9.685 220.485 -9.355 ;
        RECT 218.795 -9.685 219.125 -9.355 ;
        RECT 217.435 -9.685 217.765 -9.355 ;
        RECT 216.075 -9.685 216.405 -9.355 ;
        RECT 214.715 -9.685 215.045 -9.355 ;
        RECT 213.355 -9.685 213.685 -9.355 ;
        RECT 211.995 -9.685 212.325 -9.355 ;
        RECT 210.635 -9.685 210.965 -9.355 ;
        RECT 209.275 -9.685 209.605 -9.355 ;
        RECT 207.915 -9.685 208.245 -9.355 ;
        RECT 206.555 -9.685 206.885 -9.355 ;
        RECT 205.195 -9.685 205.525 -9.355 ;
        RECT 203.835 -9.685 204.165 -9.355 ;
        RECT 202.475 -9.685 202.805 -9.355 ;
        RECT 201.115 -9.685 201.445 -9.355 ;
        RECT 199.755 -9.685 200.085 -9.355 ;
        RECT 198.395 -9.685 198.725 -9.355 ;
        RECT 197.035 -9.685 197.365 -9.355 ;
        RECT 195.675 -9.685 196.005 -9.355 ;
        RECT 194.315 -9.685 194.645 -9.355 ;
        RECT 192.955 -9.685 193.285 -9.355 ;
        RECT 191.595 -9.685 191.925 -9.355 ;
        RECT 190.235 -9.685 190.565 -9.355 ;
        RECT 188.875 -9.685 189.205 -9.355 ;
        RECT 187.515 -9.685 187.845 -9.355 ;
        RECT 186.155 -9.685 186.485 -9.355 ;
        RECT 184.795 -9.685 185.125 -9.355 ;
        RECT 183.435 -9.685 183.765 -9.355 ;
        RECT 182.075 -9.685 182.405 -9.355 ;
        RECT 180.715 -9.685 181.045 -9.355 ;
        RECT 179.355 -9.685 179.685 -9.355 ;
        RECT 177.995 -9.685 178.325 -9.355 ;
        RECT 176.635 -9.685 176.965 -9.355 ;
        RECT 175.275 -9.685 175.605 -9.355 ;
        RECT 173.915 -9.685 174.245 -9.355 ;
        RECT 172.555 -9.685 172.885 -9.355 ;
        RECT 171.195 -9.685 171.525 -9.355 ;
        RECT 169.835 -9.685 170.165 -9.355 ;
        RECT 168.475 -9.685 168.805 -9.355 ;
        RECT 167.115 -9.685 167.445 -9.355 ;
        RECT 165.755 -9.685 166.085 -9.355 ;
        RECT 164.395 -9.685 164.725 -9.355 ;
        RECT 163.035 -9.685 163.365 -9.355 ;
        RECT 161.675 -9.685 162.005 -9.355 ;
        RECT 160.315 -9.685 160.645 -9.355 ;
        RECT 158.955 -9.685 159.285 -9.355 ;
        RECT 157.595 -9.685 157.925 -9.355 ;
        RECT 156.235 -9.685 156.565 -9.355 ;
        RECT 154.875 -9.685 155.205 -9.355 ;
        RECT 153.515 -9.685 153.845 -9.355 ;
        RECT 152.155 -9.685 152.485 -9.355 ;
        RECT 150.795 -9.685 151.125 -9.355 ;
        RECT 149.435 -9.685 149.765 -9.355 ;
        RECT 148.075 -9.685 148.405 -9.355 ;
        RECT 146.715 -9.685 147.045 -9.355 ;
        RECT 145.355 -9.685 145.685 -9.355 ;
        RECT 143.995 -9.685 144.325 -9.355 ;
        RECT 142.635 -9.685 142.965 -9.355 ;
        RECT 141.275 -9.685 141.605 -9.355 ;
        RECT 139.915 -9.685 140.245 -9.355 ;
        RECT 138.555 -9.685 138.885 -9.355 ;
        RECT 137.195 -9.685 137.525 -9.355 ;
        RECT 135.835 -9.685 136.165 -9.355 ;
        RECT 134.475 -9.685 134.805 -9.355 ;
        RECT 133.115 -9.685 133.445 -9.355 ;
        RECT 131.755 -9.685 132.085 -9.355 ;
        RECT 130.395 -9.685 130.725 -9.355 ;
        RECT 129.035 -9.685 129.365 -9.355 ;
        RECT 127.675 -9.685 128.005 -9.355 ;
        RECT 126.315 -9.685 126.645 -9.355 ;
        RECT 124.955 -9.685 125.285 -9.355 ;
        RECT 123.595 -9.685 123.925 -9.355 ;
        RECT 122.235 -9.685 122.565 -9.355 ;
        RECT 120.875 -9.685 121.205 -9.355 ;
        RECT 119.515 -9.685 119.845 -9.355 ;
        RECT 118.155 -9.685 118.485 -9.355 ;
        RECT 116.795 -9.685 117.125 -9.355 ;
        RECT 115.435 -9.685 115.765 -9.355 ;
        RECT 114.075 -9.685 114.405 -9.355 ;
        RECT 112.715 -9.685 113.045 -9.355 ;
        RECT 111.355 -9.685 111.685 -9.355 ;
        RECT 109.995 -9.685 110.325 -9.355 ;
        RECT 108.635 -9.685 108.965 -9.355 ;
        RECT 107.275 -9.685 107.605 -9.355 ;
        RECT 105.915 -9.685 106.245 -9.355 ;
        RECT 104.555 -9.685 104.885 -9.355 ;
        RECT 103.195 -9.685 103.525 -9.355 ;
        RECT 101.835 -9.685 102.165 -9.355 ;
        RECT 100.475 -9.685 100.805 -9.355 ;
        RECT 99.115 -9.685 99.445 -9.355 ;
        RECT 97.755 -9.685 98.085 -9.355 ;
        RECT 96.395 -9.685 96.725 -9.355 ;
        RECT 95.035 -9.685 95.365 -9.355 ;
        RECT 93.675 -9.685 94.005 -9.355 ;
        RECT 92.315 -9.685 92.645 -9.355 ;
        RECT 90.955 -9.685 91.285 -9.355 ;
        RECT 89.595 -9.685 89.925 -9.355 ;
        RECT 88.235 -9.685 88.565 -9.355 ;
        RECT 86.875 -9.685 87.205 -9.355 ;
        RECT 85.515 -9.685 85.845 -9.355 ;
        RECT 84.155 -9.685 84.485 -9.355 ;
        RECT 82.795 -9.685 83.125 -9.355 ;
        RECT 81.435 -9.685 81.765 -9.355 ;
        RECT 80.075 -9.685 80.405 -9.355 ;
        RECT 78.715 -9.685 79.045 -9.355 ;
        RECT 77.355 -9.685 77.685 -9.355 ;
        RECT 75.995 -9.685 76.325 -9.355 ;
        RECT 74.635 -9.685 74.965 -9.355 ;
        RECT 73.275 -9.685 73.605 -9.355 ;
        RECT 71.915 -9.685 72.245 -9.355 ;
        RECT 70.555 -9.685 70.885 -9.355 ;
        RECT 69.195 -9.685 69.525 -9.355 ;
        RECT 67.835 -9.685 68.165 -9.355 ;
        RECT 66.475 -9.685 66.805 -9.355 ;
        RECT 65.115 -9.685 65.445 -9.355 ;
        RECT 63.755 -9.685 64.085 -9.355 ;
        RECT 62.395 -9.685 62.725 -9.355 ;
        RECT 61.035 -9.685 61.365 -9.355 ;
        RECT 59.675 -9.685 60.005 -9.355 ;
        RECT 58.315 -9.685 58.645 -9.355 ;
        RECT 56.955 -9.685 57.285 -9.355 ;
        RECT 55.595 -9.685 55.925 -9.355 ;
        RECT 54.235 -9.685 54.565 -9.355 ;
        RECT 52.875 -9.685 53.205 -9.355 ;
        RECT 51.515 -9.685 51.845 -9.355 ;
        RECT 50.155 -9.685 50.485 -9.355 ;
        RECT 48.795 -9.685 49.125 -9.355 ;
        RECT 47.435 -9.685 47.765 -9.355 ;
        RECT 46.075 -9.685 46.405 -9.355 ;
        RECT 44.715 -9.685 45.045 -9.355 ;
        RECT 43.355 -9.685 43.685 -9.355 ;
        RECT 41.995 -9.685 42.325 -9.355 ;
        RECT 40.635 -9.685 40.965 -9.355 ;
        RECT 39.275 -9.685 39.605 -9.355 ;
        RECT 37.915 -9.685 38.245 -9.355 ;
        RECT 36.555 -9.685 36.885 -9.355 ;
        RECT 35.195 -9.685 35.525 -9.355 ;
        RECT 33.835 -9.685 34.165 -9.355 ;
        RECT 32.475 -9.685 32.805 -9.355 ;
        RECT 31.115 -9.685 31.445 -9.355 ;
        RECT 29.755 -9.685 30.085 -9.355 ;
        RECT 28.395 -9.685 28.725 -9.355 ;
        RECT 27.035 -9.685 27.365 -9.355 ;
        RECT 25.675 -9.685 26.005 -9.355 ;
        RECT 24.315 -9.685 24.645 -9.355 ;
        RECT 22.955 -9.685 23.285 -9.355 ;
        RECT 21.595 -9.685 21.925 -9.355 ;
        RECT 20.235 -9.685 20.565 -9.355 ;
        RECT 18.875 -9.685 19.205 -9.355 ;
        RECT 17.515 -9.685 17.845 -9.355 ;
        RECT 16.155 -9.685 16.485 -9.355 ;
        RECT 14.795 -9.685 15.125 -9.355 ;
        RECT 13.435 -9.685 13.765 -9.355 ;
        RECT 12.075 -9.685 12.405 -9.355 ;
        RECT 10.715 -9.685 11.045 -9.355 ;
        RECT 9.355 -9.685 9.685 -9.355 ;
        RECT 7.995 -9.685 8.325 -9.355 ;
        RECT 6.635 -9.685 6.965 -9.355 ;
        RECT 5.275 -9.685 5.605 -9.355 ;
        RECT 3.915 -9.685 4.245 -9.355 ;
        RECT 2.555 -9.685 2.885 -9.355 ;
        RECT 1.195 -9.685 1.525 -9.355 ;
        RECT -0.165 -9.685 0.165 -9.355 ;
        RECT -1.525 -9.685 -1.195 -9.355 ;
        RECT 954.555 -9.685 954.885 -9.355 ;
        RECT 678.475 -9.68 954.885 -9.36 ;
        RECT 953.195 -9.685 953.525 -9.355 ;
        RECT 951.835 -9.685 952.165 -9.355 ;
        RECT 950.475 -9.685 950.805 -9.355 ;
        RECT 949.115 -9.685 949.445 -9.355 ;
        RECT 947.755 -9.685 948.085 -9.355 ;
        RECT 946.395 -9.685 946.725 -9.355 ;
        RECT 945.035 -9.685 945.365 -9.355 ;
        RECT 943.675 -9.685 944.005 -9.355 ;
        RECT 942.315 -9.685 942.645 -9.355 ;
        RECT 940.955 -9.685 941.285 -9.355 ;
        RECT 939.595 -9.685 939.925 -9.355 ;
        RECT 938.235 -9.685 938.565 -9.355 ;
        RECT 936.875 -9.685 937.205 -9.355 ;
        RECT 935.515 -9.685 935.845 -9.355 ;
        RECT 934.155 -9.685 934.485 -9.355 ;
        RECT 932.795 -9.685 933.125 -9.355 ;
        RECT 931.435 -9.685 931.765 -9.355 ;
        RECT 930.075 -9.685 930.405 -9.355 ;
        RECT 928.715 -9.685 929.045 -9.355 ;
        RECT 927.355 -9.685 927.685 -9.355 ;
        RECT 925.995 -9.685 926.325 -9.355 ;
        RECT 924.635 -9.685 924.965 -9.355 ;
        RECT 923.275 -9.685 923.605 -9.355 ;
        RECT 921.915 -9.685 922.245 -9.355 ;
        RECT 920.555 -9.685 920.885 -9.355 ;
        RECT 919.195 -9.685 919.525 -9.355 ;
        RECT 917.835 -9.685 918.165 -9.355 ;
        RECT 916.475 -9.685 916.805 -9.355 ;
        RECT 915.115 -9.685 915.445 -9.355 ;
        RECT 913.755 -9.685 914.085 -9.355 ;
        RECT 912.395 -9.685 912.725 -9.355 ;
        RECT 911.035 -9.685 911.365 -9.355 ;
        RECT 909.675 -9.685 910.005 -9.355 ;
        RECT 908.315 -9.685 908.645 -9.355 ;
        RECT 906.955 -9.685 907.285 -9.355 ;
        RECT 905.595 -9.685 905.925 -9.355 ;
        RECT 904.235 -9.685 904.565 -9.355 ;
        RECT 902.875 -9.685 903.205 -9.355 ;
        RECT 901.515 -9.685 901.845 -9.355 ;
        RECT 900.155 -9.685 900.485 -9.355 ;
        RECT 898.795 -9.685 899.125 -9.355 ;
        RECT 897.435 -9.685 897.765 -9.355 ;
        RECT 896.075 -9.685 896.405 -9.355 ;
        RECT 894.715 -9.685 895.045 -9.355 ;
        RECT 893.355 -9.685 893.685 -9.355 ;
        RECT 891.995 -9.685 892.325 -9.355 ;
        RECT 890.635 -9.685 890.965 -9.355 ;
        RECT 889.275 -9.685 889.605 -9.355 ;
        RECT 887.915 -9.685 888.245 -9.355 ;
        RECT 886.555 -9.685 886.885 -9.355 ;
        RECT 885.195 -9.685 885.525 -9.355 ;
        RECT 883.835 -9.685 884.165 -9.355 ;
        RECT 882.475 -9.685 882.805 -9.355 ;
        RECT 881.115 -9.685 881.445 -9.355 ;
        RECT 879.755 -9.685 880.085 -9.355 ;
        RECT 878.395 -9.685 878.725 -9.355 ;
        RECT 877.035 -9.685 877.365 -9.355 ;
        RECT 875.675 -9.685 876.005 -9.355 ;
        RECT 874.315 -9.685 874.645 -9.355 ;
        RECT 872.955 -9.685 873.285 -9.355 ;
        RECT 871.595 -9.685 871.925 -9.355 ;
        RECT 870.235 -9.685 870.565 -9.355 ;
        RECT 868.875 -9.685 869.205 -9.355 ;
        RECT 867.515 -9.685 867.845 -9.355 ;
        RECT 866.155 -9.685 866.485 -9.355 ;
        RECT 864.795 -9.685 865.125 -9.355 ;
        RECT 863.435 -9.685 863.765 -9.355 ;
        RECT 862.075 -9.685 862.405 -9.355 ;
        RECT 860.715 -9.685 861.045 -9.355 ;
        RECT 859.355 -9.685 859.685 -9.355 ;
        RECT 857.995 -9.685 858.325 -9.355 ;
        RECT 856.635 -9.685 856.965 -9.355 ;
        RECT 855.275 -9.685 855.605 -9.355 ;
        RECT 853.915 -9.685 854.245 -9.355 ;
        RECT 852.555 -9.685 852.885 -9.355 ;
        RECT 851.195 -9.685 851.525 -9.355 ;
        RECT 849.835 -9.685 850.165 -9.355 ;
        RECT 848.475 -9.685 848.805 -9.355 ;
        RECT 847.115 -9.685 847.445 -9.355 ;
        RECT 845.755 -9.685 846.085 -9.355 ;
        RECT 844.395 -9.685 844.725 -9.355 ;
        RECT 843.035 -9.685 843.365 -9.355 ;
        RECT 841.675 -9.685 842.005 -9.355 ;
        RECT 840.315 -9.685 840.645 -9.355 ;
        RECT 838.955 -9.685 839.285 -9.355 ;
        RECT 837.595 -9.685 837.925 -9.355 ;
        RECT 836.235 -9.685 836.565 -9.355 ;
        RECT 834.875 -9.685 835.205 -9.355 ;
        RECT 833.515 -9.685 833.845 -9.355 ;
        RECT 832.155 -9.685 832.485 -9.355 ;
        RECT 830.795 -9.685 831.125 -9.355 ;
        RECT 829.435 -9.685 829.765 -9.355 ;
        RECT 828.075 -9.685 828.405 -9.355 ;
        RECT 826.715 -9.685 827.045 -9.355 ;
        RECT 825.355 -9.685 825.685 -9.355 ;
        RECT 823.995 -9.685 824.325 -9.355 ;
        RECT 822.635 -9.685 822.965 -9.355 ;
        RECT 821.275 -9.685 821.605 -9.355 ;
        RECT 819.915 -9.685 820.245 -9.355 ;
        RECT 818.555 -9.685 818.885 -9.355 ;
        RECT 817.195 -9.685 817.525 -9.355 ;
        RECT 815.835 -9.685 816.165 -9.355 ;
        RECT 814.475 -9.685 814.805 -9.355 ;
        RECT 813.115 -9.685 813.445 -9.355 ;
        RECT 811.755 -9.685 812.085 -9.355 ;
        RECT 810.395 -9.685 810.725 -9.355 ;
        RECT 809.035 -9.685 809.365 -9.355 ;
        RECT 807.675 -9.685 808.005 -9.355 ;
        RECT 806.315 -9.685 806.645 -9.355 ;
        RECT 804.955 -9.685 805.285 -9.355 ;
        RECT 803.595 -9.685 803.925 -9.355 ;
        RECT 802.235 -9.685 802.565 -9.355 ;
        RECT 800.875 -9.685 801.205 -9.355 ;
        RECT 799.515 -9.685 799.845 -9.355 ;
        RECT 798.155 -9.685 798.485 -9.355 ;
        RECT 796.795 -9.685 797.125 -9.355 ;
        RECT 795.435 -9.685 795.765 -9.355 ;
        RECT 794.075 -9.685 794.405 -9.355 ;
        RECT 792.715 -9.685 793.045 -9.355 ;
        RECT 791.355 -9.685 791.685 -9.355 ;
        RECT 789.995 -9.685 790.325 -9.355 ;
        RECT 788.635 -9.685 788.965 -9.355 ;
        RECT 787.275 -9.685 787.605 -9.355 ;
        RECT 785.915 -9.685 786.245 -9.355 ;
        RECT 784.555 -9.685 784.885 -9.355 ;
        RECT 783.195 -9.685 783.525 -9.355 ;
        RECT 781.835 -9.685 782.165 -9.355 ;
        RECT 780.475 -9.685 780.805 -9.355 ;
        RECT 779.115 -9.685 779.445 -9.355 ;
        RECT 777.755 -9.685 778.085 -9.355 ;
        RECT 776.395 -9.685 776.725 -9.355 ;
        RECT 775.035 -9.685 775.365 -9.355 ;
        RECT 773.675 -9.685 774.005 -9.355 ;
        RECT 772.315 -9.685 772.645 -9.355 ;
        RECT 770.955 -9.685 771.285 -9.355 ;
        RECT 769.595 -9.685 769.925 -9.355 ;
        RECT 768.235 -9.685 768.565 -9.355 ;
        RECT 766.875 -9.685 767.205 -9.355 ;
        RECT 765.515 -9.685 765.845 -9.355 ;
        RECT 764.155 -9.685 764.485 -9.355 ;
        RECT 762.795 -9.685 763.125 -9.355 ;
        RECT 761.435 -9.685 761.765 -9.355 ;
        RECT 760.075 -9.685 760.405 -9.355 ;
        RECT 758.715 -9.685 759.045 -9.355 ;
        RECT 757.355 -9.685 757.685 -9.355 ;
        RECT 755.995 -9.685 756.325 -9.355 ;
        RECT 754.635 -9.685 754.965 -9.355 ;
        RECT 753.275 -9.685 753.605 -9.355 ;
        RECT 751.915 -9.685 752.245 -9.355 ;
        RECT 750.555 -9.685 750.885 -9.355 ;
        RECT 749.195 -9.685 749.525 -9.355 ;
        RECT 747.835 -9.685 748.165 -9.355 ;
        RECT 746.475 -9.685 746.805 -9.355 ;
        RECT 745.115 -9.685 745.445 -9.355 ;
        RECT 743.755 -9.685 744.085 -9.355 ;
        RECT 742.395 -9.685 742.725 -9.355 ;
        RECT 741.035 -9.685 741.365 -9.355 ;
        RECT 739.675 -9.685 740.005 -9.355 ;
        RECT 738.315 -9.685 738.645 -9.355 ;
        RECT 736.955 -9.685 737.285 -9.355 ;
        RECT 735.595 -9.685 735.925 -9.355 ;
        RECT 734.235 -9.685 734.565 -9.355 ;
        RECT 732.875 -9.685 733.205 -9.355 ;
        RECT 731.515 -9.685 731.845 -9.355 ;
        RECT 730.155 -9.685 730.485 -9.355 ;
        RECT 728.795 -9.685 729.125 -9.355 ;
        RECT 727.435 -9.685 727.765 -9.355 ;
        RECT 726.075 -9.685 726.405 -9.355 ;
        RECT 724.715 -9.685 725.045 -9.355 ;
        RECT 723.355 -9.685 723.685 -9.355 ;
        RECT 721.995 -9.685 722.325 -9.355 ;
        RECT 720.635 -9.685 720.965 -9.355 ;
        RECT 719.275 -9.685 719.605 -9.355 ;
        RECT 717.915 -9.685 718.245 -9.355 ;
        RECT 716.555 -9.685 716.885 -9.355 ;
        RECT 715.195 -9.685 715.525 -9.355 ;
        RECT 713.835 -9.685 714.165 -9.355 ;
        RECT 712.475 -9.685 712.805 -9.355 ;
        RECT 711.115 -9.685 711.445 -9.355 ;
        RECT 709.755 -9.685 710.085 -9.355 ;
        RECT 708.395 -9.685 708.725 -9.355 ;
        RECT 707.035 -9.685 707.365 -9.355 ;
        RECT 705.675 -9.685 706.005 -9.355 ;
        RECT 704.315 -9.685 704.645 -9.355 ;
        RECT 702.955 -9.685 703.285 -9.355 ;
        RECT 701.595 -9.685 701.925 -9.355 ;
        RECT 700.235 -9.685 700.565 -9.355 ;
        RECT 698.875 -9.685 699.205 -9.355 ;
        RECT 697.515 -9.685 697.845 -9.355 ;
        RECT 696.155 -9.685 696.485 -9.355 ;
        RECT 694.795 -9.685 695.125 -9.355 ;
        RECT 693.435 -9.685 693.765 -9.355 ;
        RECT 692.075 -9.685 692.405 -9.355 ;
        RECT 690.715 -9.685 691.045 -9.355 ;
        RECT 689.355 -9.685 689.685 -9.355 ;
        RECT 687.995 -9.685 688.325 -9.355 ;
        RECT 686.635 -9.685 686.965 -9.355 ;
        RECT 685.275 -9.685 685.605 -9.355 ;
        RECT 683.915 -9.685 684.245 -9.355 ;
        RECT 682.555 -9.685 682.885 -9.355 ;
        RECT 681.195 -9.685 681.525 -9.355 ;
        RECT 679.835 -9.685 680.165 -9.355 ;
        RECT 678.475 -9.685 678.805 -9.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 648.555 -11.045 648.885 -10.715 ;
        RECT 647.195 -11.045 647.525 -10.715 ;
        RECT 645.835 -11.045 646.165 -10.715 ;
        RECT 644.475 -11.045 644.805 -10.715 ;
        RECT 643.115 -11.045 643.445 -10.715 ;
        RECT 641.755 -11.045 642.085 -10.715 ;
        RECT 640.395 -11.045 640.725 -10.715 ;
        RECT 639.035 -11.045 639.365 -10.715 ;
        RECT 637.675 -11.045 638.005 -10.715 ;
        RECT 636.315 -11.045 636.645 -10.715 ;
        RECT 634.955 -11.045 635.285 -10.715 ;
        RECT 633.595 -11.045 633.925 -10.715 ;
        RECT 632.235 -11.045 632.565 -10.715 ;
        RECT 630.875 -11.045 631.205 -10.715 ;
        RECT 629.515 -11.045 629.845 -10.715 ;
        RECT 628.155 -11.045 628.485 -10.715 ;
        RECT 626.795 -11.045 627.125 -10.715 ;
        RECT 625.435 -11.045 625.765 -10.715 ;
        RECT 624.075 -11.045 624.405 -10.715 ;
        RECT 622.715 -11.045 623.045 -10.715 ;
        RECT 621.355 -11.045 621.685 -10.715 ;
        RECT 619.995 -11.045 620.325 -10.715 ;
        RECT 618.635 -11.045 618.965 -10.715 ;
        RECT 617.275 -11.045 617.605 -10.715 ;
        RECT 615.915 -11.045 616.245 -10.715 ;
        RECT 614.555 -11.045 614.885 -10.715 ;
        RECT 613.195 -11.045 613.525 -10.715 ;
        RECT 611.835 -11.045 612.165 -10.715 ;
        RECT 610.475 -11.045 610.805 -10.715 ;
        RECT 609.115 -11.045 609.445 -10.715 ;
        RECT 607.755 -11.045 608.085 -10.715 ;
        RECT 606.395 -11.045 606.725 -10.715 ;
        RECT 605.035 -11.045 605.365 -10.715 ;
        RECT 603.675 -11.045 604.005 -10.715 ;
        RECT 602.315 -11.045 602.645 -10.715 ;
        RECT 600.955 -11.045 601.285 -10.715 ;
        RECT 599.595 -11.045 599.925 -10.715 ;
        RECT 598.235 -11.045 598.565 -10.715 ;
        RECT 596.875 -11.045 597.205 -10.715 ;
        RECT 595.515 -11.045 595.845 -10.715 ;
        RECT 594.155 -11.045 594.485 -10.715 ;
        RECT 592.795 -11.045 593.125 -10.715 ;
        RECT 591.435 -11.045 591.765 -10.715 ;
        RECT 590.075 -11.045 590.405 -10.715 ;
        RECT 588.715 -11.045 589.045 -10.715 ;
        RECT 587.355 -11.045 587.685 -10.715 ;
        RECT 585.995 -11.045 586.325 -10.715 ;
        RECT 584.635 -11.045 584.965 -10.715 ;
        RECT 583.275 -11.045 583.605 -10.715 ;
        RECT 581.915 -11.045 582.245 -10.715 ;
        RECT 580.555 -11.045 580.885 -10.715 ;
        RECT 579.195 -11.045 579.525 -10.715 ;
        RECT 577.835 -11.045 578.165 -10.715 ;
        RECT 576.475 -11.045 576.805 -10.715 ;
        RECT 575.115 -11.045 575.445 -10.715 ;
        RECT 573.755 -11.045 574.085 -10.715 ;
        RECT 572.395 -11.045 572.725 -10.715 ;
        RECT 571.035 -11.045 571.365 -10.715 ;
        RECT 569.675 -11.045 570.005 -10.715 ;
        RECT 568.315 -11.045 568.645 -10.715 ;
        RECT 566.955 -11.045 567.285 -10.715 ;
        RECT 565.595 -11.045 565.925 -10.715 ;
        RECT 564.235 -11.045 564.565 -10.715 ;
        RECT 562.875 -11.045 563.205 -10.715 ;
        RECT 561.515 -11.045 561.845 -10.715 ;
        RECT 560.155 -11.045 560.485 -10.715 ;
        RECT 558.795 -11.045 559.125 -10.715 ;
        RECT 557.435 -11.045 557.765 -10.715 ;
        RECT 556.075 -11.045 556.405 -10.715 ;
        RECT 554.715 -11.045 555.045 -10.715 ;
        RECT 553.355 -11.045 553.685 -10.715 ;
        RECT 551.995 -11.045 552.325 -10.715 ;
        RECT 550.635 -11.045 550.965 -10.715 ;
        RECT 549.275 -11.045 549.605 -10.715 ;
        RECT 547.915 -11.045 548.245 -10.715 ;
        RECT 546.555 -11.045 546.885 -10.715 ;
        RECT 545.195 -11.045 545.525 -10.715 ;
        RECT 543.835 -11.045 544.165 -10.715 ;
        RECT 542.475 -11.045 542.805 -10.715 ;
        RECT 541.115 -11.045 541.445 -10.715 ;
        RECT 539.755 -11.045 540.085 -10.715 ;
        RECT 538.395 -11.045 538.725 -10.715 ;
        RECT 537.035 -11.045 537.365 -10.715 ;
        RECT 535.675 -11.045 536.005 -10.715 ;
        RECT 534.315 -11.045 534.645 -10.715 ;
        RECT 532.955 -11.045 533.285 -10.715 ;
        RECT 531.595 -11.045 531.925 -10.715 ;
        RECT 530.235 -11.045 530.565 -10.715 ;
        RECT 528.875 -11.045 529.205 -10.715 ;
        RECT 527.515 -11.045 527.845 -10.715 ;
        RECT 526.155 -11.045 526.485 -10.715 ;
        RECT 524.795 -11.045 525.125 -10.715 ;
        RECT 523.435 -11.045 523.765 -10.715 ;
        RECT 522.075 -11.045 522.405 -10.715 ;
        RECT 520.715 -11.045 521.045 -10.715 ;
        RECT 519.355 -11.045 519.685 -10.715 ;
        RECT 517.995 -11.045 518.325 -10.715 ;
        RECT 516.635 -11.045 516.965 -10.715 ;
        RECT 515.275 -11.045 515.605 -10.715 ;
        RECT 513.915 -11.045 514.245 -10.715 ;
        RECT 512.555 -11.045 512.885 -10.715 ;
        RECT 511.195 -11.045 511.525 -10.715 ;
        RECT 509.835 -11.045 510.165 -10.715 ;
        RECT 508.475 -11.045 508.805 -10.715 ;
        RECT 507.115 -11.045 507.445 -10.715 ;
        RECT 505.755 -11.045 506.085 -10.715 ;
        RECT 504.395 -11.045 504.725 -10.715 ;
        RECT 503.035 -11.045 503.365 -10.715 ;
        RECT 501.675 -11.045 502.005 -10.715 ;
        RECT 500.315 -11.045 500.645 -10.715 ;
        RECT 498.955 -11.045 499.285 -10.715 ;
        RECT 497.595 -11.045 497.925 -10.715 ;
        RECT 496.235 -11.045 496.565 -10.715 ;
        RECT 494.875 -11.045 495.205 -10.715 ;
        RECT 493.515 -11.045 493.845 -10.715 ;
        RECT 492.155 -11.045 492.485 -10.715 ;
        RECT 490.795 -11.045 491.125 -10.715 ;
        RECT 489.435 -11.045 489.765 -10.715 ;
        RECT 488.075 -11.045 488.405 -10.715 ;
        RECT 486.715 -11.045 487.045 -10.715 ;
        RECT 485.355 -11.045 485.685 -10.715 ;
        RECT 483.995 -11.045 484.325 -10.715 ;
        RECT 482.635 -11.045 482.965 -10.715 ;
        RECT 481.275 -11.045 481.605 -10.715 ;
        RECT 479.915 -11.045 480.245 -10.715 ;
        RECT 478.555 -11.045 478.885 -10.715 ;
        RECT 477.195 -11.045 477.525 -10.715 ;
        RECT 475.835 -11.045 476.165 -10.715 ;
        RECT 474.475 -11.045 474.805 -10.715 ;
        RECT 473.115 -11.045 473.445 -10.715 ;
        RECT 471.755 -11.045 472.085 -10.715 ;
        RECT 470.395 -11.045 470.725 -10.715 ;
        RECT 469.035 -11.045 469.365 -10.715 ;
        RECT 467.675 -11.045 468.005 -10.715 ;
        RECT 466.315 -11.045 466.645 -10.715 ;
        RECT 464.955 -11.045 465.285 -10.715 ;
        RECT 463.595 -11.045 463.925 -10.715 ;
        RECT 462.235 -11.045 462.565 -10.715 ;
        RECT 460.875 -11.045 461.205 -10.715 ;
        RECT 459.515 -11.045 459.845 -10.715 ;
        RECT 458.155 -11.045 458.485 -10.715 ;
        RECT 456.795 -11.045 457.125 -10.715 ;
        RECT 455.435 -11.045 455.765 -10.715 ;
        RECT 454.075 -11.045 454.405 -10.715 ;
        RECT 452.715 -11.045 453.045 -10.715 ;
        RECT 451.355 -11.045 451.685 -10.715 ;
        RECT 449.995 -11.045 450.325 -10.715 ;
        RECT 448.635 -11.045 448.965 -10.715 ;
        RECT 447.275 -11.045 447.605 -10.715 ;
        RECT 445.915 -11.045 446.245 -10.715 ;
        RECT 444.555 -11.045 444.885 -10.715 ;
        RECT 443.195 -11.045 443.525 -10.715 ;
        RECT 441.835 -11.045 442.165 -10.715 ;
        RECT 440.475 -11.045 440.805 -10.715 ;
        RECT 439.115 -11.045 439.445 -10.715 ;
        RECT 437.755 -11.045 438.085 -10.715 ;
        RECT 436.395 -11.045 436.725 -10.715 ;
        RECT 435.035 -11.045 435.365 -10.715 ;
        RECT 433.675 -11.045 434.005 -10.715 ;
        RECT 432.315 -11.045 432.645 -10.715 ;
        RECT 430.955 -11.045 431.285 -10.715 ;
        RECT 429.595 -11.045 429.925 -10.715 ;
        RECT 428.235 -11.045 428.565 -10.715 ;
        RECT 426.875 -11.045 427.205 -10.715 ;
        RECT 425.515 -11.045 425.845 -10.715 ;
        RECT 424.155 -11.045 424.485 -10.715 ;
        RECT 422.795 -11.045 423.125 -10.715 ;
        RECT 421.435 -11.045 421.765 -10.715 ;
        RECT 420.075 -11.045 420.405 -10.715 ;
        RECT 418.715 -11.045 419.045 -10.715 ;
        RECT 417.355 -11.045 417.685 -10.715 ;
        RECT 415.995 -11.045 416.325 -10.715 ;
        RECT 414.635 -11.045 414.965 -10.715 ;
        RECT 413.275 -11.045 413.605 -10.715 ;
        RECT 411.915 -11.045 412.245 -10.715 ;
        RECT 410.555 -11.045 410.885 -10.715 ;
        RECT 409.195 -11.045 409.525 -10.715 ;
        RECT 407.835 -11.045 408.165 -10.715 ;
        RECT 406.475 -11.045 406.805 -10.715 ;
        RECT 405.115 -11.045 405.445 -10.715 ;
        RECT 403.755 -11.045 404.085 -10.715 ;
        RECT 402.395 -11.045 402.725 -10.715 ;
        RECT 401.035 -11.045 401.365 -10.715 ;
        RECT 399.675 -11.045 400.005 -10.715 ;
        RECT 398.315 -11.045 398.645 -10.715 ;
        RECT 396.955 -11.045 397.285 -10.715 ;
        RECT 395.595 -11.045 395.925 -10.715 ;
        RECT 394.235 -11.045 394.565 -10.715 ;
        RECT 392.875 -11.045 393.205 -10.715 ;
        RECT 391.515 -11.045 391.845 -10.715 ;
        RECT 390.155 -11.045 390.485 -10.715 ;
        RECT 388.795 -11.045 389.125 -10.715 ;
        RECT 387.435 -11.045 387.765 -10.715 ;
        RECT 386.075 -11.045 386.405 -10.715 ;
        RECT 384.715 -11.045 385.045 -10.715 ;
        RECT 383.355 -11.045 383.685 -10.715 ;
        RECT 381.995 -11.045 382.325 -10.715 ;
        RECT 380.635 -11.045 380.965 -10.715 ;
        RECT 379.275 -11.045 379.605 -10.715 ;
        RECT 377.915 -11.045 378.245 -10.715 ;
        RECT 376.555 -11.045 376.885 -10.715 ;
        RECT 375.195 -11.045 375.525 -10.715 ;
        RECT 373.835 -11.045 374.165 -10.715 ;
        RECT 372.475 -11.045 372.805 -10.715 ;
        RECT 371.115 -11.045 371.445 -10.715 ;
        RECT 369.755 -11.045 370.085 -10.715 ;
        RECT 368.395 -11.045 368.725 -10.715 ;
        RECT 367.035 -11.045 367.365 -10.715 ;
        RECT 365.675 -11.045 366.005 -10.715 ;
        RECT 364.315 -11.045 364.645 -10.715 ;
        RECT 362.955 -11.045 363.285 -10.715 ;
        RECT 361.595 -11.045 361.925 -10.715 ;
        RECT 360.235 -11.045 360.565 -10.715 ;
        RECT 358.875 -11.045 359.205 -10.715 ;
        RECT 357.515 -11.045 357.845 -10.715 ;
        RECT 356.155 -11.045 356.485 -10.715 ;
        RECT 354.795 -11.045 355.125 -10.715 ;
        RECT 353.435 -11.045 353.765 -10.715 ;
        RECT 352.075 -11.045 352.405 -10.715 ;
        RECT 350.715 -11.045 351.045 -10.715 ;
        RECT 349.355 -11.045 349.685 -10.715 ;
        RECT 347.995 -11.045 348.325 -10.715 ;
        RECT 346.635 -11.045 346.965 -10.715 ;
        RECT 345.275 -11.045 345.605 -10.715 ;
        RECT 343.915 -11.045 344.245 -10.715 ;
        RECT 342.555 -11.045 342.885 -10.715 ;
        RECT 341.195 -11.045 341.525 -10.715 ;
        RECT 339.835 -11.045 340.165 -10.715 ;
        RECT 338.475 -11.045 338.805 -10.715 ;
        RECT 337.115 -11.045 337.445 -10.715 ;
        RECT 335.755 -11.045 336.085 -10.715 ;
        RECT 334.395 -11.045 334.725 -10.715 ;
        RECT 333.035 -11.045 333.365 -10.715 ;
        RECT 331.675 -11.045 332.005 -10.715 ;
        RECT 330.315 -11.045 330.645 -10.715 ;
        RECT 328.955 -11.045 329.285 -10.715 ;
        RECT 327.595 -11.045 327.925 -10.715 ;
        RECT 326.235 -11.045 326.565 -10.715 ;
        RECT 324.875 -11.045 325.205 -10.715 ;
        RECT 323.515 -11.045 323.845 -10.715 ;
        RECT 322.155 -11.045 322.485 -10.715 ;
        RECT 320.795 -11.045 321.125 -10.715 ;
        RECT 319.435 -11.045 319.765 -10.715 ;
        RECT 318.075 -11.045 318.405 -10.715 ;
        RECT 316.715 -11.045 317.045 -10.715 ;
        RECT 315.355 -11.045 315.685 -10.715 ;
        RECT 313.995 -11.045 314.325 -10.715 ;
        RECT 312.635 -11.045 312.965 -10.715 ;
        RECT 311.275 -11.045 311.605 -10.715 ;
        RECT 309.915 -11.045 310.245 -10.715 ;
        RECT 308.555 -11.045 308.885 -10.715 ;
        RECT 307.195 -11.045 307.525 -10.715 ;
        RECT 305.835 -11.045 306.165 -10.715 ;
        RECT 304.475 -11.045 304.805 -10.715 ;
        RECT 303.115 -11.045 303.445 -10.715 ;
        RECT 301.755 -11.045 302.085 -10.715 ;
        RECT 300.395 -11.045 300.725 -10.715 ;
        RECT 299.035 -11.045 299.365 -10.715 ;
        RECT 297.675 -11.045 298.005 -10.715 ;
        RECT 296.315 -11.045 296.645 -10.715 ;
        RECT 294.955 -11.045 295.285 -10.715 ;
        RECT 293.595 -11.045 293.925 -10.715 ;
        RECT 292.235 -11.045 292.565 -10.715 ;
        RECT 290.875 -11.045 291.205 -10.715 ;
        RECT 289.515 -11.045 289.845 -10.715 ;
        RECT 288.155 -11.045 288.485 -10.715 ;
        RECT 286.795 -11.045 287.125 -10.715 ;
        RECT 285.435 -11.045 285.765 -10.715 ;
        RECT 284.075 -11.045 284.405 -10.715 ;
        RECT 282.715 -11.045 283.045 -10.715 ;
        RECT 281.355 -11.045 281.685 -10.715 ;
        RECT 279.995 -11.045 280.325 -10.715 ;
        RECT 278.635 -11.045 278.965 -10.715 ;
        RECT 277.275 -11.045 277.605 -10.715 ;
        RECT 275.915 -11.045 276.245 -10.715 ;
        RECT 274.555 -11.045 274.885 -10.715 ;
        RECT 273.195 -11.045 273.525 -10.715 ;
        RECT 271.835 -11.045 272.165 -10.715 ;
        RECT 270.475 -11.045 270.805 -10.715 ;
        RECT 269.115 -11.045 269.445 -10.715 ;
        RECT 267.755 -11.045 268.085 -10.715 ;
        RECT 266.395 -11.045 266.725 -10.715 ;
        RECT 265.035 -11.045 265.365 -10.715 ;
        RECT 263.675 -11.045 264.005 -10.715 ;
        RECT 262.315 -11.045 262.645 -10.715 ;
        RECT 260.955 -11.045 261.285 -10.715 ;
        RECT 259.595 -11.045 259.925 -10.715 ;
        RECT 258.235 -11.045 258.565 -10.715 ;
        RECT 256.875 -11.045 257.205 -10.715 ;
        RECT 255.515 -11.045 255.845 -10.715 ;
        RECT 254.155 -11.045 254.485 -10.715 ;
        RECT 252.795 -11.045 253.125 -10.715 ;
        RECT 251.435 -11.045 251.765 -10.715 ;
        RECT 250.075 -11.045 250.405 -10.715 ;
        RECT 248.715 -11.045 249.045 -10.715 ;
        RECT 247.355 -11.045 247.685 -10.715 ;
        RECT 245.995 -11.045 246.325 -10.715 ;
        RECT 244.635 -11.045 244.965 -10.715 ;
        RECT 243.275 -11.045 243.605 -10.715 ;
        RECT 241.915 -11.045 242.245 -10.715 ;
        RECT 240.555 -11.045 240.885 -10.715 ;
        RECT 239.195 -11.045 239.525 -10.715 ;
        RECT 237.835 -11.045 238.165 -10.715 ;
        RECT 236.475 -11.045 236.805 -10.715 ;
        RECT 235.115 -11.045 235.445 -10.715 ;
        RECT 233.755 -11.045 234.085 -10.715 ;
        RECT 232.395 -11.045 232.725 -10.715 ;
        RECT 231.035 -11.045 231.365 -10.715 ;
        RECT 229.675 -11.045 230.005 -10.715 ;
        RECT 228.315 -11.045 228.645 -10.715 ;
        RECT 226.955 -11.045 227.285 -10.715 ;
        RECT 225.595 -11.045 225.925 -10.715 ;
        RECT 224.235 -11.045 224.565 -10.715 ;
        RECT 222.875 -11.045 223.205 -10.715 ;
        RECT 221.515 -11.045 221.845 -10.715 ;
        RECT 220.155 -11.045 220.485 -10.715 ;
        RECT 218.795 -11.045 219.125 -10.715 ;
        RECT 217.435 -11.045 217.765 -10.715 ;
        RECT 216.075 -11.045 216.405 -10.715 ;
        RECT 214.715 -11.045 215.045 -10.715 ;
        RECT 213.355 -11.045 213.685 -10.715 ;
        RECT 211.995 -11.045 212.325 -10.715 ;
        RECT 210.635 -11.045 210.965 -10.715 ;
        RECT 209.275 -11.045 209.605 -10.715 ;
        RECT 207.915 -11.045 208.245 -10.715 ;
        RECT 206.555 -11.045 206.885 -10.715 ;
        RECT 205.195 -11.045 205.525 -10.715 ;
        RECT 203.835 -11.045 204.165 -10.715 ;
        RECT 202.475 -11.045 202.805 -10.715 ;
        RECT 201.115 -11.045 201.445 -10.715 ;
        RECT 199.755 -11.045 200.085 -10.715 ;
        RECT 198.395 -11.045 198.725 -10.715 ;
        RECT 197.035 -11.045 197.365 -10.715 ;
        RECT 195.675 -11.045 196.005 -10.715 ;
        RECT 194.315 -11.045 194.645 -10.715 ;
        RECT 192.955 -11.045 193.285 -10.715 ;
        RECT 191.595 -11.045 191.925 -10.715 ;
        RECT 190.235 -11.045 190.565 -10.715 ;
        RECT 188.875 -11.045 189.205 -10.715 ;
        RECT 187.515 -11.045 187.845 -10.715 ;
        RECT 186.155 -11.045 186.485 -10.715 ;
        RECT 184.795 -11.045 185.125 -10.715 ;
        RECT 183.435 -11.045 183.765 -10.715 ;
        RECT 182.075 -11.045 182.405 -10.715 ;
        RECT 180.715 -11.045 181.045 -10.715 ;
        RECT 179.355 -11.045 179.685 -10.715 ;
        RECT 177.995 -11.045 178.325 -10.715 ;
        RECT 176.635 -11.045 176.965 -10.715 ;
        RECT 175.275 -11.045 175.605 -10.715 ;
        RECT 173.915 -11.045 174.245 -10.715 ;
        RECT 172.555 -11.045 172.885 -10.715 ;
        RECT 171.195 -11.045 171.525 -10.715 ;
        RECT 169.835 -11.045 170.165 -10.715 ;
        RECT 168.475 -11.045 168.805 -10.715 ;
        RECT 167.115 -11.045 167.445 -10.715 ;
        RECT 165.755 -11.045 166.085 -10.715 ;
        RECT 164.395 -11.045 164.725 -10.715 ;
        RECT 163.035 -11.045 163.365 -10.715 ;
        RECT 161.675 -11.045 162.005 -10.715 ;
        RECT 160.315 -11.045 160.645 -10.715 ;
        RECT 158.955 -11.045 159.285 -10.715 ;
        RECT 157.595 -11.045 157.925 -10.715 ;
        RECT 156.235 -11.045 156.565 -10.715 ;
        RECT 154.875 -11.045 155.205 -10.715 ;
        RECT 153.515 -11.045 153.845 -10.715 ;
        RECT 152.155 -11.045 152.485 -10.715 ;
        RECT 150.795 -11.045 151.125 -10.715 ;
        RECT 149.435 -11.045 149.765 -10.715 ;
        RECT 148.075 -11.045 148.405 -10.715 ;
        RECT 146.715 -11.045 147.045 -10.715 ;
        RECT 145.355 -11.045 145.685 -10.715 ;
        RECT 143.995 -11.045 144.325 -10.715 ;
        RECT 142.635 -11.045 142.965 -10.715 ;
        RECT 141.275 -11.045 141.605 -10.715 ;
        RECT 139.915 -11.045 140.245 -10.715 ;
        RECT 138.555 -11.045 138.885 -10.715 ;
        RECT 137.195 -11.045 137.525 -10.715 ;
        RECT 135.835 -11.045 136.165 -10.715 ;
        RECT 134.475 -11.045 134.805 -10.715 ;
        RECT 133.115 -11.045 133.445 -10.715 ;
        RECT 131.755 -11.045 132.085 -10.715 ;
        RECT 130.395 -11.045 130.725 -10.715 ;
        RECT 129.035 -11.045 129.365 -10.715 ;
        RECT 127.675 -11.045 128.005 -10.715 ;
        RECT 126.315 -11.045 126.645 -10.715 ;
        RECT 124.955 -11.045 125.285 -10.715 ;
        RECT 123.595 -11.045 123.925 -10.715 ;
        RECT 122.235 -11.045 122.565 -10.715 ;
        RECT 120.875 -11.045 121.205 -10.715 ;
        RECT 119.515 -11.045 119.845 -10.715 ;
        RECT 118.155 -11.045 118.485 -10.715 ;
        RECT 116.795 -11.045 117.125 -10.715 ;
        RECT 115.435 -11.045 115.765 -10.715 ;
        RECT 114.075 -11.045 114.405 -10.715 ;
        RECT 112.715 -11.045 113.045 -10.715 ;
        RECT 111.355 -11.045 111.685 -10.715 ;
        RECT 109.995 -11.045 110.325 -10.715 ;
        RECT 108.635 -11.045 108.965 -10.715 ;
        RECT 107.275 -11.045 107.605 -10.715 ;
        RECT 105.915 -11.045 106.245 -10.715 ;
        RECT 104.555 -11.045 104.885 -10.715 ;
        RECT 103.195 -11.045 103.525 -10.715 ;
        RECT 101.835 -11.045 102.165 -10.715 ;
        RECT 100.475 -11.045 100.805 -10.715 ;
        RECT 99.115 -11.045 99.445 -10.715 ;
        RECT 97.755 -11.045 98.085 -10.715 ;
        RECT 96.395 -11.045 96.725 -10.715 ;
        RECT 95.035 -11.045 95.365 -10.715 ;
        RECT 93.675 -11.045 94.005 -10.715 ;
        RECT 92.315 -11.045 92.645 -10.715 ;
        RECT 90.955 -11.045 91.285 -10.715 ;
        RECT 89.595 -11.045 89.925 -10.715 ;
        RECT 88.235 -11.045 88.565 -10.715 ;
        RECT 86.875 -11.045 87.205 -10.715 ;
        RECT 85.515 -11.045 85.845 -10.715 ;
        RECT 84.155 -11.045 84.485 -10.715 ;
        RECT 82.795 -11.045 83.125 -10.715 ;
        RECT 81.435 -11.045 81.765 -10.715 ;
        RECT 80.075 -11.045 80.405 -10.715 ;
        RECT 78.715 -11.045 79.045 -10.715 ;
        RECT 77.355 -11.045 77.685 -10.715 ;
        RECT 75.995 -11.045 76.325 -10.715 ;
        RECT 74.635 -11.045 74.965 -10.715 ;
        RECT 73.275 -11.045 73.605 -10.715 ;
        RECT 71.915 -11.045 72.245 -10.715 ;
        RECT 70.555 -11.045 70.885 -10.715 ;
        RECT 69.195 -11.045 69.525 -10.715 ;
        RECT 67.835 -11.045 68.165 -10.715 ;
        RECT 66.475 -11.045 66.805 -10.715 ;
        RECT 65.115 -11.045 65.445 -10.715 ;
        RECT 63.755 -11.045 64.085 -10.715 ;
        RECT 62.395 -11.045 62.725 -10.715 ;
        RECT 61.035 -11.045 61.365 -10.715 ;
        RECT 59.675 -11.045 60.005 -10.715 ;
        RECT 58.315 -11.045 58.645 -10.715 ;
        RECT 56.955 -11.045 57.285 -10.715 ;
        RECT 55.595 -11.045 55.925 -10.715 ;
        RECT 54.235 -11.045 54.565 -10.715 ;
        RECT 52.875 -11.045 53.205 -10.715 ;
        RECT 51.515 -11.045 51.845 -10.715 ;
        RECT 50.155 -11.045 50.485 -10.715 ;
        RECT 48.795 -11.045 49.125 -10.715 ;
        RECT 47.435 -11.045 47.765 -10.715 ;
        RECT 46.075 -11.045 46.405 -10.715 ;
        RECT 44.715 -11.045 45.045 -10.715 ;
        RECT 43.355 -11.045 43.685 -10.715 ;
        RECT 41.995 -11.045 42.325 -10.715 ;
        RECT 40.635 -11.045 40.965 -10.715 ;
        RECT 39.275 -11.045 39.605 -10.715 ;
        RECT 37.915 -11.045 38.245 -10.715 ;
        RECT 36.555 -11.045 36.885 -10.715 ;
        RECT 35.195 -11.045 35.525 -10.715 ;
        RECT 33.835 -11.045 34.165 -10.715 ;
        RECT 32.475 -11.045 32.805 -10.715 ;
        RECT 31.115 -11.045 31.445 -10.715 ;
        RECT 29.755 -11.045 30.085 -10.715 ;
        RECT 28.395 -11.045 28.725 -10.715 ;
        RECT 27.035 -11.045 27.365 -10.715 ;
        RECT 25.675 -11.045 26.005 -10.715 ;
        RECT 24.315 -11.045 24.645 -10.715 ;
        RECT 22.955 -11.045 23.285 -10.715 ;
        RECT 21.595 -11.045 21.925 -10.715 ;
        RECT 20.235 -11.045 20.565 -10.715 ;
        RECT 18.875 -11.045 19.205 -10.715 ;
        RECT 17.515 -11.045 17.845 -10.715 ;
        RECT 16.155 -11.045 16.485 -10.715 ;
        RECT 14.795 -11.045 15.125 -10.715 ;
        RECT 13.435 -11.045 13.765 -10.715 ;
        RECT 12.075 -11.045 12.405 -10.715 ;
        RECT 10.715 -11.045 11.045 -10.715 ;
        RECT 9.355 -11.045 9.685 -10.715 ;
        RECT 7.995 -11.045 8.325 -10.715 ;
        RECT 6.635 -11.045 6.965 -10.715 ;
        RECT 5.275 -11.045 5.605 -10.715 ;
        RECT 3.915 -11.045 4.245 -10.715 ;
        RECT 2.555 -11.045 2.885 -10.715 ;
        RECT 1.195 -11.045 1.525 -10.715 ;
        RECT -0.165 -11.045 0.165 -10.715 ;
        RECT -1.525 -11.045 -1.195 -10.715 ;
        RECT -1.525 -11.04 678.475 -10.72 ;
        RECT 677.115 -11.045 677.445 -10.715 ;
        RECT 675.755 -11.045 676.085 -10.715 ;
        RECT 674.395 -11.045 674.725 -10.715 ;
        RECT 673.035 -11.045 673.365 -10.715 ;
        RECT 671.675 -11.045 672.005 -10.715 ;
        RECT 670.315 -11.045 670.645 -10.715 ;
        RECT 668.955 -11.045 669.285 -10.715 ;
        RECT 667.595 -11.045 667.925 -10.715 ;
        RECT 666.235 -11.045 666.565 -10.715 ;
        RECT 664.875 -11.045 665.205 -10.715 ;
        RECT 663.515 -11.045 663.845 -10.715 ;
        RECT 662.155 -11.045 662.485 -10.715 ;
        RECT 660.795 -11.045 661.125 -10.715 ;
        RECT 659.435 -11.045 659.765 -10.715 ;
        RECT 658.075 -11.045 658.405 -10.715 ;
        RECT 656.715 -11.045 657.045 -10.715 ;
        RECT 655.355 -11.045 655.685 -10.715 ;
        RECT 653.995 -11.045 654.325 -10.715 ;
        RECT 652.635 -11.045 652.965 -10.715 ;
        RECT 651.275 -11.045 651.605 -10.715 ;
        RECT 649.915 -11.045 650.245 -10.715 ;
        RECT 840.315 -11.045 840.645 -10.715 ;
        RECT 838.955 -11.045 839.285 -10.715 ;
        RECT 837.595 -11.045 837.925 -10.715 ;
        RECT 836.235 -11.045 836.565 -10.715 ;
        RECT 834.875 -11.045 835.205 -10.715 ;
        RECT 833.515 -11.045 833.845 -10.715 ;
        RECT 832.155 -11.045 832.485 -10.715 ;
        RECT 830.795 -11.045 831.125 -10.715 ;
        RECT 829.435 -11.045 829.765 -10.715 ;
        RECT 828.075 -11.045 828.405 -10.715 ;
        RECT 826.715 -11.045 827.045 -10.715 ;
        RECT 825.355 -11.045 825.685 -10.715 ;
        RECT 823.995 -11.045 824.325 -10.715 ;
        RECT 822.635 -11.045 822.965 -10.715 ;
        RECT 821.275 -11.045 821.605 -10.715 ;
        RECT 819.915 -11.045 820.245 -10.715 ;
        RECT 818.555 -11.045 818.885 -10.715 ;
        RECT 817.195 -11.045 817.525 -10.715 ;
        RECT 815.835 -11.045 816.165 -10.715 ;
        RECT 814.475 -11.045 814.805 -10.715 ;
        RECT 813.115 -11.045 813.445 -10.715 ;
        RECT 811.755 -11.045 812.085 -10.715 ;
        RECT 810.395 -11.045 810.725 -10.715 ;
        RECT 809.035 -11.045 809.365 -10.715 ;
        RECT 807.675 -11.045 808.005 -10.715 ;
        RECT 806.315 -11.045 806.645 -10.715 ;
        RECT 804.955 -11.045 805.285 -10.715 ;
        RECT 803.595 -11.045 803.925 -10.715 ;
        RECT 802.235 -11.045 802.565 -10.715 ;
        RECT 800.875 -11.045 801.205 -10.715 ;
        RECT 799.515 -11.045 799.845 -10.715 ;
        RECT 798.155 -11.045 798.485 -10.715 ;
        RECT 796.795 -11.045 797.125 -10.715 ;
        RECT 795.435 -11.045 795.765 -10.715 ;
        RECT 794.075 -11.045 794.405 -10.715 ;
        RECT 792.715 -11.045 793.045 -10.715 ;
        RECT 791.355 -11.045 791.685 -10.715 ;
        RECT 789.995 -11.045 790.325 -10.715 ;
        RECT 788.635 -11.045 788.965 -10.715 ;
        RECT 787.275 -11.045 787.605 -10.715 ;
        RECT 785.915 -11.045 786.245 -10.715 ;
        RECT 784.555 -11.045 784.885 -10.715 ;
        RECT 783.195 -11.045 783.525 -10.715 ;
        RECT 781.835 -11.045 782.165 -10.715 ;
        RECT 780.475 -11.045 780.805 -10.715 ;
        RECT 779.115 -11.045 779.445 -10.715 ;
        RECT 777.755 -11.045 778.085 -10.715 ;
        RECT 776.395 -11.045 776.725 -10.715 ;
        RECT 775.035 -11.045 775.365 -10.715 ;
        RECT 773.675 -11.045 774.005 -10.715 ;
        RECT 772.315 -11.045 772.645 -10.715 ;
        RECT 770.955 -11.045 771.285 -10.715 ;
        RECT 769.595 -11.045 769.925 -10.715 ;
        RECT 768.235 -11.045 768.565 -10.715 ;
        RECT 766.875 -11.045 767.205 -10.715 ;
        RECT 765.515 -11.045 765.845 -10.715 ;
        RECT 764.155 -11.045 764.485 -10.715 ;
        RECT 762.795 -11.045 763.125 -10.715 ;
        RECT 761.435 -11.045 761.765 -10.715 ;
        RECT 760.075 -11.045 760.405 -10.715 ;
        RECT 758.715 -11.045 759.045 -10.715 ;
        RECT 757.355 -11.045 757.685 -10.715 ;
        RECT 755.995 -11.045 756.325 -10.715 ;
        RECT 754.635 -11.045 754.965 -10.715 ;
        RECT 753.275 -11.045 753.605 -10.715 ;
        RECT 751.915 -11.045 752.245 -10.715 ;
        RECT 750.555 -11.045 750.885 -10.715 ;
        RECT 749.195 -11.045 749.525 -10.715 ;
        RECT 747.835 -11.045 748.165 -10.715 ;
        RECT 746.475 -11.045 746.805 -10.715 ;
        RECT 745.115 -11.045 745.445 -10.715 ;
        RECT 743.755 -11.045 744.085 -10.715 ;
        RECT 742.395 -11.045 742.725 -10.715 ;
        RECT 741.035 -11.045 741.365 -10.715 ;
        RECT 739.675 -11.045 740.005 -10.715 ;
        RECT 738.315 -11.045 738.645 -10.715 ;
        RECT 736.955 -11.045 737.285 -10.715 ;
        RECT 735.595 -11.045 735.925 -10.715 ;
        RECT 734.235 -11.045 734.565 -10.715 ;
        RECT 732.875 -11.045 733.205 -10.715 ;
        RECT 731.515 -11.045 731.845 -10.715 ;
        RECT 730.155 -11.045 730.485 -10.715 ;
        RECT 728.795 -11.045 729.125 -10.715 ;
        RECT 727.435 -11.045 727.765 -10.715 ;
        RECT 726.075 -11.045 726.405 -10.715 ;
        RECT 724.715 -11.045 725.045 -10.715 ;
        RECT 723.355 -11.045 723.685 -10.715 ;
        RECT 721.995 -11.045 722.325 -10.715 ;
        RECT 720.635 -11.045 720.965 -10.715 ;
        RECT 719.275 -11.045 719.605 -10.715 ;
        RECT 717.915 -11.045 718.245 -10.715 ;
        RECT 716.555 -11.045 716.885 -10.715 ;
        RECT 715.195 -11.045 715.525 -10.715 ;
        RECT 713.835 -11.045 714.165 -10.715 ;
        RECT 712.475 -11.045 712.805 -10.715 ;
        RECT 711.115 -11.045 711.445 -10.715 ;
        RECT 709.755 -11.045 710.085 -10.715 ;
        RECT 708.395 -11.045 708.725 -10.715 ;
        RECT 707.035 -11.045 707.365 -10.715 ;
        RECT 705.675 -11.045 706.005 -10.715 ;
        RECT 704.315 -11.045 704.645 -10.715 ;
        RECT 702.955 -11.045 703.285 -10.715 ;
        RECT 701.595 -11.045 701.925 -10.715 ;
        RECT 700.235 -11.045 700.565 -10.715 ;
        RECT 698.875 -11.045 699.205 -10.715 ;
        RECT 697.515 -11.045 697.845 -10.715 ;
        RECT 696.155 -11.045 696.485 -10.715 ;
        RECT 694.795 -11.045 695.125 -10.715 ;
        RECT 693.435 -11.045 693.765 -10.715 ;
        RECT 692.075 -11.045 692.405 -10.715 ;
        RECT 690.715 -11.045 691.045 -10.715 ;
        RECT 689.355 -11.045 689.685 -10.715 ;
        RECT 687.995 -11.045 688.325 -10.715 ;
        RECT 686.635 -11.045 686.965 -10.715 ;
        RECT 685.275 -11.045 685.605 -10.715 ;
        RECT 683.915 -11.045 684.245 -10.715 ;
        RECT 682.555 -11.045 682.885 -10.715 ;
        RECT 681.195 -11.045 681.525 -10.715 ;
        RECT 679.835 -11.045 680.165 -10.715 ;
        RECT 678.475 -11.045 678.805 -10.715 ;
        RECT 954.555 -11.045 954.885 -10.715 ;
        RECT 678.475 -11.04 954.885 -10.72 ;
        RECT 953.195 -11.045 953.525 -10.715 ;
        RECT 951.835 -11.045 952.165 -10.715 ;
        RECT 950.475 -11.045 950.805 -10.715 ;
        RECT 949.115 -11.045 949.445 -10.715 ;
        RECT 947.755 -11.045 948.085 -10.715 ;
        RECT 946.395 -11.045 946.725 -10.715 ;
        RECT 945.035 -11.045 945.365 -10.715 ;
        RECT 943.675 -11.045 944.005 -10.715 ;
        RECT 942.315 -11.045 942.645 -10.715 ;
        RECT 940.955 -11.045 941.285 -10.715 ;
        RECT 939.595 -11.045 939.925 -10.715 ;
        RECT 938.235 -11.045 938.565 -10.715 ;
        RECT 936.875 -11.045 937.205 -10.715 ;
        RECT 935.515 -11.045 935.845 -10.715 ;
        RECT 934.155 -11.045 934.485 -10.715 ;
        RECT 932.795 -11.045 933.125 -10.715 ;
        RECT 931.435 -11.045 931.765 -10.715 ;
        RECT 930.075 -11.045 930.405 -10.715 ;
        RECT 928.715 -11.045 929.045 -10.715 ;
        RECT 927.355 -11.045 927.685 -10.715 ;
        RECT 925.995 -11.045 926.325 -10.715 ;
        RECT 924.635 -11.045 924.965 -10.715 ;
        RECT 923.275 -11.045 923.605 -10.715 ;
        RECT 921.915 -11.045 922.245 -10.715 ;
        RECT 920.555 -11.045 920.885 -10.715 ;
        RECT 919.195 -11.045 919.525 -10.715 ;
        RECT 917.835 -11.045 918.165 -10.715 ;
        RECT 916.475 -11.045 916.805 -10.715 ;
        RECT 915.115 -11.045 915.445 -10.715 ;
        RECT 913.755 -11.045 914.085 -10.715 ;
        RECT 912.395 -11.045 912.725 -10.715 ;
        RECT 911.035 -11.045 911.365 -10.715 ;
        RECT 909.675 -11.045 910.005 -10.715 ;
        RECT 908.315 -11.045 908.645 -10.715 ;
        RECT 906.955 -11.045 907.285 -10.715 ;
        RECT 905.595 -11.045 905.925 -10.715 ;
        RECT 904.235 -11.045 904.565 -10.715 ;
        RECT 902.875 -11.045 903.205 -10.715 ;
        RECT 901.515 -11.045 901.845 -10.715 ;
        RECT 900.155 -11.045 900.485 -10.715 ;
        RECT 898.795 -11.045 899.125 -10.715 ;
        RECT 897.435 -11.045 897.765 -10.715 ;
        RECT 896.075 -11.045 896.405 -10.715 ;
        RECT 894.715 -11.045 895.045 -10.715 ;
        RECT 893.355 -11.045 893.685 -10.715 ;
        RECT 891.995 -11.045 892.325 -10.715 ;
        RECT 890.635 -11.045 890.965 -10.715 ;
        RECT 889.275 -11.045 889.605 -10.715 ;
        RECT 887.915 -11.045 888.245 -10.715 ;
        RECT 886.555 -11.045 886.885 -10.715 ;
        RECT 885.195 -11.045 885.525 -10.715 ;
        RECT 883.835 -11.045 884.165 -10.715 ;
        RECT 882.475 -11.045 882.805 -10.715 ;
        RECT 881.115 -11.045 881.445 -10.715 ;
        RECT 879.755 -11.045 880.085 -10.715 ;
        RECT 878.395 -11.045 878.725 -10.715 ;
        RECT 877.035 -11.045 877.365 -10.715 ;
        RECT 875.675 -11.045 876.005 -10.715 ;
        RECT 874.315 -11.045 874.645 -10.715 ;
        RECT 872.955 -11.045 873.285 -10.715 ;
        RECT 871.595 -11.045 871.925 -10.715 ;
        RECT 870.235 -11.045 870.565 -10.715 ;
        RECT 868.875 -11.045 869.205 -10.715 ;
        RECT 867.515 -11.045 867.845 -10.715 ;
        RECT 866.155 -11.045 866.485 -10.715 ;
        RECT 864.795 -11.045 865.125 -10.715 ;
        RECT 863.435 -11.045 863.765 -10.715 ;
        RECT 862.075 -11.045 862.405 -10.715 ;
        RECT 860.715 -11.045 861.045 -10.715 ;
        RECT 859.355 -11.045 859.685 -10.715 ;
        RECT 857.995 -11.045 858.325 -10.715 ;
        RECT 856.635 -11.045 856.965 -10.715 ;
        RECT 855.275 -11.045 855.605 -10.715 ;
        RECT 853.915 -11.045 854.245 -10.715 ;
        RECT 852.555 -11.045 852.885 -10.715 ;
        RECT 851.195 -11.045 851.525 -10.715 ;
        RECT 849.835 -11.045 850.165 -10.715 ;
        RECT 848.475 -11.045 848.805 -10.715 ;
        RECT 847.115 -11.045 847.445 -10.715 ;
        RECT 845.755 -11.045 846.085 -10.715 ;
        RECT 844.395 -11.045 844.725 -10.715 ;
        RECT 843.035 -11.045 843.365 -10.715 ;
        RECT 841.675 -11.045 842.005 -10.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -6.96 678.475 -6.64 ;
        RECT 677.115 -6.965 677.445 -6.635 ;
        RECT 675.755 -6.965 676.085 -6.635 ;
        RECT 674.395 -6.965 674.725 -6.635 ;
        RECT 673.035 -6.965 673.365 -6.635 ;
        RECT 671.675 -6.965 672.005 -6.635 ;
        RECT 670.315 -6.965 670.645 -6.635 ;
        RECT 668.955 -6.965 669.285 -6.635 ;
        RECT 667.595 -6.965 667.925 -6.635 ;
        RECT 666.235 -6.965 666.565 -6.635 ;
        RECT 664.875 -6.965 665.205 -6.635 ;
        RECT 663.515 -6.965 663.845 -6.635 ;
        RECT 662.155 -6.965 662.485 -6.635 ;
        RECT 660.795 -6.965 661.125 -6.635 ;
        RECT 659.435 -6.965 659.765 -6.635 ;
        RECT 658.075 -6.965 658.405 -6.635 ;
        RECT 656.715 -6.965 657.045 -6.635 ;
        RECT 655.355 -6.965 655.685 -6.635 ;
        RECT 653.995 -6.965 654.325 -6.635 ;
        RECT 652.635 -6.965 652.965 -6.635 ;
        RECT 651.275 -6.965 651.605 -6.635 ;
        RECT 649.915 -6.965 650.245 -6.635 ;
        RECT 648.555 -6.965 648.885 -6.635 ;
        RECT 647.195 -6.965 647.525 -6.635 ;
        RECT 645.835 -6.965 646.165 -6.635 ;
        RECT 644.475 -6.965 644.805 -6.635 ;
        RECT 643.115 -6.965 643.445 -6.635 ;
        RECT 641.755 -6.965 642.085 -6.635 ;
        RECT 640.395 -6.965 640.725 -6.635 ;
        RECT 639.035 -6.965 639.365 -6.635 ;
        RECT 637.675 -6.965 638.005 -6.635 ;
        RECT 636.315 -6.965 636.645 -6.635 ;
        RECT 634.955 -6.965 635.285 -6.635 ;
        RECT 633.595 -6.965 633.925 -6.635 ;
        RECT 632.235 -6.965 632.565 -6.635 ;
        RECT 630.875 -6.965 631.205 -6.635 ;
        RECT 629.515 -6.965 629.845 -6.635 ;
        RECT 628.155 -6.965 628.485 -6.635 ;
        RECT 626.795 -6.965 627.125 -6.635 ;
        RECT 625.435 -6.965 625.765 -6.635 ;
        RECT 624.075 -6.965 624.405 -6.635 ;
        RECT 622.715 -6.965 623.045 -6.635 ;
        RECT 621.355 -6.965 621.685 -6.635 ;
        RECT 619.995 -6.965 620.325 -6.635 ;
        RECT 618.635 -6.965 618.965 -6.635 ;
        RECT 617.275 -6.965 617.605 -6.635 ;
        RECT 615.915 -6.965 616.245 -6.635 ;
        RECT 614.555 -6.965 614.885 -6.635 ;
        RECT 613.195 -6.965 613.525 -6.635 ;
        RECT 611.835 -6.965 612.165 -6.635 ;
        RECT 610.475 -6.965 610.805 -6.635 ;
        RECT 609.115 -6.965 609.445 -6.635 ;
        RECT 607.755 -6.965 608.085 -6.635 ;
        RECT 606.395 -6.965 606.725 -6.635 ;
        RECT 605.035 -6.965 605.365 -6.635 ;
        RECT 603.675 -6.965 604.005 -6.635 ;
        RECT 602.315 -6.965 602.645 -6.635 ;
        RECT 600.955 -6.965 601.285 -6.635 ;
        RECT 599.595 -6.965 599.925 -6.635 ;
        RECT 598.235 -6.965 598.565 -6.635 ;
        RECT 596.875 -6.965 597.205 -6.635 ;
        RECT 595.515 -6.965 595.845 -6.635 ;
        RECT 594.155 -6.965 594.485 -6.635 ;
        RECT 592.795 -6.965 593.125 -6.635 ;
        RECT 591.435 -6.965 591.765 -6.635 ;
        RECT 590.075 -6.965 590.405 -6.635 ;
        RECT 588.715 -6.965 589.045 -6.635 ;
        RECT 587.355 -6.965 587.685 -6.635 ;
        RECT 585.995 -6.965 586.325 -6.635 ;
        RECT 584.635 -6.965 584.965 -6.635 ;
        RECT 583.275 -6.965 583.605 -6.635 ;
        RECT 581.915 -6.965 582.245 -6.635 ;
        RECT 580.555 -6.965 580.885 -6.635 ;
        RECT 579.195 -6.965 579.525 -6.635 ;
        RECT 577.835 -6.965 578.165 -6.635 ;
        RECT 576.475 -6.965 576.805 -6.635 ;
        RECT 575.115 -6.965 575.445 -6.635 ;
        RECT 573.755 -6.965 574.085 -6.635 ;
        RECT 572.395 -6.965 572.725 -6.635 ;
        RECT 571.035 -6.965 571.365 -6.635 ;
        RECT 569.675 -6.965 570.005 -6.635 ;
        RECT 568.315 -6.965 568.645 -6.635 ;
        RECT 566.955 -6.965 567.285 -6.635 ;
        RECT 565.595 -6.965 565.925 -6.635 ;
        RECT 564.235 -6.965 564.565 -6.635 ;
        RECT 562.875 -6.965 563.205 -6.635 ;
        RECT 561.515 -6.965 561.845 -6.635 ;
        RECT 560.155 -6.965 560.485 -6.635 ;
        RECT 558.795 -6.965 559.125 -6.635 ;
        RECT 557.435 -6.965 557.765 -6.635 ;
        RECT 556.075 -6.965 556.405 -6.635 ;
        RECT 554.715 -6.965 555.045 -6.635 ;
        RECT 553.355 -6.965 553.685 -6.635 ;
        RECT 551.995 -6.965 552.325 -6.635 ;
        RECT 550.635 -6.965 550.965 -6.635 ;
        RECT 549.275 -6.965 549.605 -6.635 ;
        RECT 547.915 -6.965 548.245 -6.635 ;
        RECT 546.555 -6.965 546.885 -6.635 ;
        RECT 545.195 -6.965 545.525 -6.635 ;
        RECT 543.835 -6.965 544.165 -6.635 ;
        RECT 542.475 -6.965 542.805 -6.635 ;
        RECT 541.115 -6.965 541.445 -6.635 ;
        RECT 539.755 -6.965 540.085 -6.635 ;
        RECT 538.395 -6.965 538.725 -6.635 ;
        RECT 537.035 -6.965 537.365 -6.635 ;
        RECT 535.675 -6.965 536.005 -6.635 ;
        RECT 534.315 -6.965 534.645 -6.635 ;
        RECT 532.955 -6.965 533.285 -6.635 ;
        RECT 531.595 -6.965 531.925 -6.635 ;
        RECT 530.235 -6.965 530.565 -6.635 ;
        RECT 528.875 -6.965 529.205 -6.635 ;
        RECT 527.515 -6.965 527.845 -6.635 ;
        RECT 526.155 -6.965 526.485 -6.635 ;
        RECT 524.795 -6.965 525.125 -6.635 ;
        RECT 523.435 -6.965 523.765 -6.635 ;
        RECT 522.075 -6.965 522.405 -6.635 ;
        RECT 520.715 -6.965 521.045 -6.635 ;
        RECT 519.355 -6.965 519.685 -6.635 ;
        RECT 517.995 -6.965 518.325 -6.635 ;
        RECT 516.635 -6.965 516.965 -6.635 ;
        RECT 515.275 -6.965 515.605 -6.635 ;
        RECT 513.915 -6.965 514.245 -6.635 ;
        RECT 512.555 -6.965 512.885 -6.635 ;
        RECT 511.195 -6.965 511.525 -6.635 ;
        RECT 509.835 -6.965 510.165 -6.635 ;
        RECT 508.475 -6.965 508.805 -6.635 ;
        RECT 507.115 -6.965 507.445 -6.635 ;
        RECT 505.755 -6.965 506.085 -6.635 ;
        RECT 504.395 -6.965 504.725 -6.635 ;
        RECT 503.035 -6.965 503.365 -6.635 ;
        RECT 501.675 -6.965 502.005 -6.635 ;
        RECT 500.315 -6.965 500.645 -6.635 ;
        RECT 498.955 -6.965 499.285 -6.635 ;
        RECT 497.595 -6.965 497.925 -6.635 ;
        RECT 496.235 -6.965 496.565 -6.635 ;
        RECT 494.875 -6.965 495.205 -6.635 ;
        RECT 493.515 -6.965 493.845 -6.635 ;
        RECT 492.155 -6.965 492.485 -6.635 ;
        RECT 490.795 -6.965 491.125 -6.635 ;
        RECT 489.435 -6.965 489.765 -6.635 ;
        RECT 488.075 -6.965 488.405 -6.635 ;
        RECT 486.715 -6.965 487.045 -6.635 ;
        RECT 485.355 -6.965 485.685 -6.635 ;
        RECT 483.995 -6.965 484.325 -6.635 ;
        RECT 482.635 -6.965 482.965 -6.635 ;
        RECT 481.275 -6.965 481.605 -6.635 ;
        RECT 479.915 -6.965 480.245 -6.635 ;
        RECT 478.555 -6.965 478.885 -6.635 ;
        RECT 477.195 -6.965 477.525 -6.635 ;
        RECT 475.835 -6.965 476.165 -6.635 ;
        RECT 474.475 -6.965 474.805 -6.635 ;
        RECT 473.115 -6.965 473.445 -6.635 ;
        RECT 471.755 -6.965 472.085 -6.635 ;
        RECT 470.395 -6.965 470.725 -6.635 ;
        RECT 469.035 -6.965 469.365 -6.635 ;
        RECT 467.675 -6.965 468.005 -6.635 ;
        RECT 466.315 -6.965 466.645 -6.635 ;
        RECT 464.955 -6.965 465.285 -6.635 ;
        RECT 463.595 -6.965 463.925 -6.635 ;
        RECT 462.235 -6.965 462.565 -6.635 ;
        RECT 460.875 -6.965 461.205 -6.635 ;
        RECT 459.515 -6.965 459.845 -6.635 ;
        RECT 458.155 -6.965 458.485 -6.635 ;
        RECT 456.795 -6.965 457.125 -6.635 ;
        RECT 455.435 -6.965 455.765 -6.635 ;
        RECT 454.075 -6.965 454.405 -6.635 ;
        RECT 452.715 -6.965 453.045 -6.635 ;
        RECT 451.355 -6.965 451.685 -6.635 ;
        RECT 449.995 -6.965 450.325 -6.635 ;
        RECT 448.635 -6.965 448.965 -6.635 ;
        RECT 447.275 -6.965 447.605 -6.635 ;
        RECT 445.915 -6.965 446.245 -6.635 ;
        RECT 444.555 -6.965 444.885 -6.635 ;
        RECT 443.195 -6.965 443.525 -6.635 ;
        RECT 441.835 -6.965 442.165 -6.635 ;
        RECT 440.475 -6.965 440.805 -6.635 ;
        RECT 439.115 -6.965 439.445 -6.635 ;
        RECT 437.755 -6.965 438.085 -6.635 ;
        RECT 436.395 -6.965 436.725 -6.635 ;
        RECT 435.035 -6.965 435.365 -6.635 ;
        RECT 433.675 -6.965 434.005 -6.635 ;
        RECT 432.315 -6.965 432.645 -6.635 ;
        RECT 430.955 -6.965 431.285 -6.635 ;
        RECT 429.595 -6.965 429.925 -6.635 ;
        RECT 428.235 -6.965 428.565 -6.635 ;
        RECT 426.875 -6.965 427.205 -6.635 ;
        RECT 425.515 -6.965 425.845 -6.635 ;
        RECT 424.155 -6.965 424.485 -6.635 ;
        RECT 422.795 -6.965 423.125 -6.635 ;
        RECT 421.435 -6.965 421.765 -6.635 ;
        RECT 420.075 -6.965 420.405 -6.635 ;
        RECT 418.715 -6.965 419.045 -6.635 ;
        RECT 417.355 -6.965 417.685 -6.635 ;
        RECT 415.995 -6.965 416.325 -6.635 ;
        RECT 414.635 -6.965 414.965 -6.635 ;
        RECT 413.275 -6.965 413.605 -6.635 ;
        RECT 411.915 -6.965 412.245 -6.635 ;
        RECT 410.555 -6.965 410.885 -6.635 ;
        RECT 409.195 -6.965 409.525 -6.635 ;
        RECT 407.835 -6.965 408.165 -6.635 ;
        RECT 406.475 -6.965 406.805 -6.635 ;
        RECT 405.115 -6.965 405.445 -6.635 ;
        RECT 403.755 -6.965 404.085 -6.635 ;
        RECT 402.395 -6.965 402.725 -6.635 ;
        RECT 401.035 -6.965 401.365 -6.635 ;
        RECT 399.675 -6.965 400.005 -6.635 ;
        RECT 398.315 -6.965 398.645 -6.635 ;
        RECT 396.955 -6.965 397.285 -6.635 ;
        RECT 395.595 -6.965 395.925 -6.635 ;
        RECT 394.235 -6.965 394.565 -6.635 ;
        RECT 392.875 -6.965 393.205 -6.635 ;
        RECT 391.515 -6.965 391.845 -6.635 ;
        RECT 390.155 -6.965 390.485 -6.635 ;
        RECT 388.795 -6.965 389.125 -6.635 ;
        RECT 387.435 -6.965 387.765 -6.635 ;
        RECT 386.075 -6.965 386.405 -6.635 ;
        RECT 384.715 -6.965 385.045 -6.635 ;
        RECT 383.355 -6.965 383.685 -6.635 ;
        RECT 381.995 -6.965 382.325 -6.635 ;
        RECT 380.635 -6.965 380.965 -6.635 ;
        RECT 379.275 -6.965 379.605 -6.635 ;
        RECT 377.915 -6.965 378.245 -6.635 ;
        RECT 376.555 -6.965 376.885 -6.635 ;
        RECT 375.195 -6.965 375.525 -6.635 ;
        RECT 373.835 -6.965 374.165 -6.635 ;
        RECT 372.475 -6.965 372.805 -6.635 ;
        RECT 371.115 -6.965 371.445 -6.635 ;
        RECT 369.755 -6.965 370.085 -6.635 ;
        RECT 368.395 -6.965 368.725 -6.635 ;
        RECT 367.035 -6.965 367.365 -6.635 ;
        RECT 365.675 -6.965 366.005 -6.635 ;
        RECT 364.315 -6.965 364.645 -6.635 ;
        RECT 362.955 -6.965 363.285 -6.635 ;
        RECT 361.595 -6.965 361.925 -6.635 ;
        RECT 360.235 -6.965 360.565 -6.635 ;
        RECT 358.875 -6.965 359.205 -6.635 ;
        RECT 357.515 -6.965 357.845 -6.635 ;
        RECT 356.155 -6.965 356.485 -6.635 ;
        RECT 354.795 -6.965 355.125 -6.635 ;
        RECT 353.435 -6.965 353.765 -6.635 ;
        RECT 352.075 -6.965 352.405 -6.635 ;
        RECT 350.715 -6.965 351.045 -6.635 ;
        RECT 349.355 -6.965 349.685 -6.635 ;
        RECT 347.995 -6.965 348.325 -6.635 ;
        RECT 346.635 -6.965 346.965 -6.635 ;
        RECT 345.275 -6.965 345.605 -6.635 ;
        RECT 343.915 -6.965 344.245 -6.635 ;
        RECT 342.555 -6.965 342.885 -6.635 ;
        RECT 341.195 -6.965 341.525 -6.635 ;
        RECT 339.835 -6.965 340.165 -6.635 ;
        RECT 338.475 -6.965 338.805 -6.635 ;
        RECT 337.115 -6.965 337.445 -6.635 ;
        RECT 335.755 -6.965 336.085 -6.635 ;
        RECT 334.395 -6.965 334.725 -6.635 ;
        RECT 333.035 -6.965 333.365 -6.635 ;
        RECT 331.675 -6.965 332.005 -6.635 ;
        RECT 330.315 -6.965 330.645 -6.635 ;
        RECT 328.955 -6.965 329.285 -6.635 ;
        RECT 327.595 -6.965 327.925 -6.635 ;
        RECT 326.235 -6.965 326.565 -6.635 ;
        RECT 324.875 -6.965 325.205 -6.635 ;
        RECT 323.515 -6.965 323.845 -6.635 ;
        RECT 322.155 -6.965 322.485 -6.635 ;
        RECT 320.795 -6.965 321.125 -6.635 ;
        RECT 319.435 -6.965 319.765 -6.635 ;
        RECT 318.075 -6.965 318.405 -6.635 ;
        RECT 316.715 -6.965 317.045 -6.635 ;
        RECT 315.355 -6.965 315.685 -6.635 ;
        RECT 313.995 -6.965 314.325 -6.635 ;
        RECT 312.635 -6.965 312.965 -6.635 ;
        RECT 311.275 -6.965 311.605 -6.635 ;
        RECT 309.915 -6.965 310.245 -6.635 ;
        RECT 308.555 -6.965 308.885 -6.635 ;
        RECT 307.195 -6.965 307.525 -6.635 ;
        RECT 305.835 -6.965 306.165 -6.635 ;
        RECT 304.475 -6.965 304.805 -6.635 ;
        RECT 303.115 -6.965 303.445 -6.635 ;
        RECT 301.755 -6.965 302.085 -6.635 ;
        RECT 300.395 -6.965 300.725 -6.635 ;
        RECT 299.035 -6.965 299.365 -6.635 ;
        RECT 297.675 -6.965 298.005 -6.635 ;
        RECT 296.315 -6.965 296.645 -6.635 ;
        RECT 294.955 -6.965 295.285 -6.635 ;
        RECT 293.595 -6.965 293.925 -6.635 ;
        RECT 292.235 -6.965 292.565 -6.635 ;
        RECT 290.875 -6.965 291.205 -6.635 ;
        RECT 289.515 -6.965 289.845 -6.635 ;
        RECT 288.155 -6.965 288.485 -6.635 ;
        RECT 286.795 -6.965 287.125 -6.635 ;
        RECT 285.435 -6.965 285.765 -6.635 ;
        RECT 284.075 -6.965 284.405 -6.635 ;
        RECT 282.715 -6.965 283.045 -6.635 ;
        RECT 281.355 -6.965 281.685 -6.635 ;
        RECT 279.995 -6.965 280.325 -6.635 ;
        RECT 278.635 -6.965 278.965 -6.635 ;
        RECT 277.275 -6.965 277.605 -6.635 ;
        RECT 275.915 -6.965 276.245 -6.635 ;
        RECT 274.555 -6.965 274.885 -6.635 ;
        RECT 273.195 -6.965 273.525 -6.635 ;
        RECT 271.835 -6.965 272.165 -6.635 ;
        RECT 270.475 -6.965 270.805 -6.635 ;
        RECT 269.115 -6.965 269.445 -6.635 ;
        RECT 267.755 -6.965 268.085 -6.635 ;
        RECT 266.395 -6.965 266.725 -6.635 ;
        RECT 265.035 -6.965 265.365 -6.635 ;
        RECT 263.675 -6.965 264.005 -6.635 ;
        RECT 262.315 -6.965 262.645 -6.635 ;
        RECT 260.955 -6.965 261.285 -6.635 ;
        RECT 259.595 -6.965 259.925 -6.635 ;
        RECT 258.235 -6.965 258.565 -6.635 ;
        RECT 256.875 -6.965 257.205 -6.635 ;
        RECT 255.515 -6.965 255.845 -6.635 ;
        RECT 254.155 -6.965 254.485 -6.635 ;
        RECT 252.795 -6.965 253.125 -6.635 ;
        RECT 251.435 -6.965 251.765 -6.635 ;
        RECT 250.075 -6.965 250.405 -6.635 ;
        RECT 248.715 -6.965 249.045 -6.635 ;
        RECT 247.355 -6.965 247.685 -6.635 ;
        RECT 245.995 -6.965 246.325 -6.635 ;
        RECT 244.635 -6.965 244.965 -6.635 ;
        RECT 243.275 -6.965 243.605 -6.635 ;
        RECT 241.915 -6.965 242.245 -6.635 ;
        RECT 240.555 -6.965 240.885 -6.635 ;
        RECT 239.195 -6.965 239.525 -6.635 ;
        RECT 237.835 -6.965 238.165 -6.635 ;
        RECT 236.475 -6.965 236.805 -6.635 ;
        RECT 235.115 -6.965 235.445 -6.635 ;
        RECT 233.755 -6.965 234.085 -6.635 ;
        RECT 232.395 -6.965 232.725 -6.635 ;
        RECT 231.035 -6.965 231.365 -6.635 ;
        RECT 229.675 -6.965 230.005 -6.635 ;
        RECT 228.315 -6.965 228.645 -6.635 ;
        RECT 226.955 -6.965 227.285 -6.635 ;
        RECT 225.595 -6.965 225.925 -6.635 ;
        RECT 224.235 -6.965 224.565 -6.635 ;
        RECT 222.875 -6.965 223.205 -6.635 ;
        RECT 221.515 -6.965 221.845 -6.635 ;
        RECT 220.155 -6.965 220.485 -6.635 ;
        RECT 218.795 -6.965 219.125 -6.635 ;
        RECT 217.435 -6.965 217.765 -6.635 ;
        RECT 216.075 -6.965 216.405 -6.635 ;
        RECT 214.715 -6.965 215.045 -6.635 ;
        RECT 213.355 -6.965 213.685 -6.635 ;
        RECT 211.995 -6.965 212.325 -6.635 ;
        RECT 210.635 -6.965 210.965 -6.635 ;
        RECT 209.275 -6.965 209.605 -6.635 ;
        RECT 207.915 -6.965 208.245 -6.635 ;
        RECT 206.555 -6.965 206.885 -6.635 ;
        RECT 205.195 -6.965 205.525 -6.635 ;
        RECT 203.835 -6.965 204.165 -6.635 ;
        RECT 202.475 -6.965 202.805 -6.635 ;
        RECT 201.115 -6.965 201.445 -6.635 ;
        RECT 199.755 -6.965 200.085 -6.635 ;
        RECT 198.395 -6.965 198.725 -6.635 ;
        RECT 197.035 -6.965 197.365 -6.635 ;
        RECT 195.675 -6.965 196.005 -6.635 ;
        RECT 194.315 -6.965 194.645 -6.635 ;
        RECT 192.955 -6.965 193.285 -6.635 ;
        RECT 191.595 -6.965 191.925 -6.635 ;
        RECT 190.235 -6.965 190.565 -6.635 ;
        RECT 188.875 -6.965 189.205 -6.635 ;
        RECT 187.515 -6.965 187.845 -6.635 ;
        RECT 186.155 -6.965 186.485 -6.635 ;
        RECT 184.795 -6.965 185.125 -6.635 ;
        RECT 183.435 -6.965 183.765 -6.635 ;
        RECT 182.075 -6.965 182.405 -6.635 ;
        RECT 180.715 -6.965 181.045 -6.635 ;
        RECT 179.355 -6.965 179.685 -6.635 ;
        RECT 177.995 -6.965 178.325 -6.635 ;
        RECT 176.635 -6.965 176.965 -6.635 ;
        RECT 175.275 -6.965 175.605 -6.635 ;
        RECT 173.915 -6.965 174.245 -6.635 ;
        RECT 172.555 -6.965 172.885 -6.635 ;
        RECT 171.195 -6.965 171.525 -6.635 ;
        RECT 169.835 -6.965 170.165 -6.635 ;
        RECT 168.475 -6.965 168.805 -6.635 ;
        RECT 167.115 -6.965 167.445 -6.635 ;
        RECT 165.755 -6.965 166.085 -6.635 ;
        RECT 164.395 -6.965 164.725 -6.635 ;
        RECT 163.035 -6.965 163.365 -6.635 ;
        RECT 161.675 -6.965 162.005 -6.635 ;
        RECT 160.315 -6.965 160.645 -6.635 ;
        RECT 158.955 -6.965 159.285 -6.635 ;
        RECT 157.595 -6.965 157.925 -6.635 ;
        RECT 156.235 -6.965 156.565 -6.635 ;
        RECT 154.875 -6.965 155.205 -6.635 ;
        RECT 153.515 -6.965 153.845 -6.635 ;
        RECT 152.155 -6.965 152.485 -6.635 ;
        RECT 150.795 -6.965 151.125 -6.635 ;
        RECT 149.435 -6.965 149.765 -6.635 ;
        RECT 148.075 -6.965 148.405 -6.635 ;
        RECT 146.715 -6.965 147.045 -6.635 ;
        RECT 145.355 -6.965 145.685 -6.635 ;
        RECT 143.995 -6.965 144.325 -6.635 ;
        RECT 142.635 -6.965 142.965 -6.635 ;
        RECT 141.275 -6.965 141.605 -6.635 ;
        RECT 139.915 -6.965 140.245 -6.635 ;
        RECT 138.555 -6.965 138.885 -6.635 ;
        RECT 137.195 -6.965 137.525 -6.635 ;
        RECT 135.835 -6.965 136.165 -6.635 ;
        RECT 134.475 -6.965 134.805 -6.635 ;
        RECT 133.115 -6.965 133.445 -6.635 ;
        RECT 131.755 -6.965 132.085 -6.635 ;
        RECT 130.395 -6.965 130.725 -6.635 ;
        RECT 129.035 -6.965 129.365 -6.635 ;
        RECT 127.675 -6.965 128.005 -6.635 ;
        RECT 126.315 -6.965 126.645 -6.635 ;
        RECT 124.955 -6.965 125.285 -6.635 ;
        RECT 123.595 -6.965 123.925 -6.635 ;
        RECT 122.235 -6.965 122.565 -6.635 ;
        RECT 120.875 -6.965 121.205 -6.635 ;
        RECT 119.515 -6.965 119.845 -6.635 ;
        RECT 118.155 -6.965 118.485 -6.635 ;
        RECT 116.795 -6.965 117.125 -6.635 ;
        RECT 115.435 -6.965 115.765 -6.635 ;
        RECT 114.075 -6.965 114.405 -6.635 ;
        RECT 112.715 -6.965 113.045 -6.635 ;
        RECT 111.355 -6.965 111.685 -6.635 ;
        RECT 109.995 -6.965 110.325 -6.635 ;
        RECT 108.635 -6.965 108.965 -6.635 ;
        RECT 107.275 -6.965 107.605 -6.635 ;
        RECT 105.915 -6.965 106.245 -6.635 ;
        RECT 104.555 -6.965 104.885 -6.635 ;
        RECT 103.195 -6.965 103.525 -6.635 ;
        RECT 101.835 -6.965 102.165 -6.635 ;
        RECT 100.475 -6.965 100.805 -6.635 ;
        RECT 99.115 -6.965 99.445 -6.635 ;
        RECT 97.755 -6.965 98.085 -6.635 ;
        RECT 96.395 -6.965 96.725 -6.635 ;
        RECT 95.035 -6.965 95.365 -6.635 ;
        RECT 93.675 -6.965 94.005 -6.635 ;
        RECT 92.315 -6.965 92.645 -6.635 ;
        RECT 90.955 -6.965 91.285 -6.635 ;
        RECT 89.595 -6.965 89.925 -6.635 ;
        RECT 88.235 -6.965 88.565 -6.635 ;
        RECT 86.875 -6.965 87.205 -6.635 ;
        RECT 85.515 -6.965 85.845 -6.635 ;
        RECT 84.155 -6.965 84.485 -6.635 ;
        RECT 82.795 -6.965 83.125 -6.635 ;
        RECT 81.435 -6.965 81.765 -6.635 ;
        RECT 80.075 -6.965 80.405 -6.635 ;
        RECT 78.715 -6.965 79.045 -6.635 ;
        RECT 77.355 -6.965 77.685 -6.635 ;
        RECT 75.995 -6.965 76.325 -6.635 ;
        RECT 74.635 -6.965 74.965 -6.635 ;
        RECT 73.275 -6.965 73.605 -6.635 ;
        RECT 71.915 -6.965 72.245 -6.635 ;
        RECT 70.555 -6.965 70.885 -6.635 ;
        RECT 69.195 -6.965 69.525 -6.635 ;
        RECT 67.835 -6.965 68.165 -6.635 ;
        RECT 66.475 -6.965 66.805 -6.635 ;
        RECT 65.115 -6.965 65.445 -6.635 ;
        RECT 63.755 -6.965 64.085 -6.635 ;
        RECT 62.395 -6.965 62.725 -6.635 ;
        RECT 61.035 -6.965 61.365 -6.635 ;
        RECT 59.675 -6.965 60.005 -6.635 ;
        RECT 58.315 -6.965 58.645 -6.635 ;
        RECT 56.955 -6.965 57.285 -6.635 ;
        RECT 55.595 -6.965 55.925 -6.635 ;
        RECT 54.235 -6.965 54.565 -6.635 ;
        RECT 52.875 -6.965 53.205 -6.635 ;
        RECT 51.515 -6.965 51.845 -6.635 ;
        RECT 50.155 -6.965 50.485 -6.635 ;
        RECT 48.795 -6.965 49.125 -6.635 ;
        RECT 47.435 -6.965 47.765 -6.635 ;
        RECT 46.075 -6.965 46.405 -6.635 ;
        RECT 44.715 -6.965 45.045 -6.635 ;
        RECT 43.355 -6.965 43.685 -6.635 ;
        RECT 41.995 -6.965 42.325 -6.635 ;
        RECT 40.635 -6.965 40.965 -6.635 ;
        RECT 39.275 -6.965 39.605 -6.635 ;
        RECT 37.915 -6.965 38.245 -6.635 ;
        RECT 36.555 -6.965 36.885 -6.635 ;
        RECT 35.195 -6.965 35.525 -6.635 ;
        RECT 33.835 -6.965 34.165 -6.635 ;
        RECT 32.475 -6.965 32.805 -6.635 ;
        RECT 31.115 -6.965 31.445 -6.635 ;
        RECT 29.755 -6.965 30.085 -6.635 ;
        RECT 28.395 -6.965 28.725 -6.635 ;
        RECT 27.035 -6.965 27.365 -6.635 ;
        RECT 25.675 -6.965 26.005 -6.635 ;
        RECT 24.315 -6.965 24.645 -6.635 ;
        RECT 22.955 -6.965 23.285 -6.635 ;
        RECT 21.595 -6.965 21.925 -6.635 ;
        RECT 20.235 -6.965 20.565 -6.635 ;
        RECT 18.875 -6.965 19.205 -6.635 ;
        RECT 17.515 -6.965 17.845 -6.635 ;
        RECT 16.155 -6.965 16.485 -6.635 ;
        RECT 14.795 -6.965 15.125 -6.635 ;
        RECT 13.435 -6.965 13.765 -6.635 ;
        RECT 12.075 -6.965 12.405 -6.635 ;
        RECT 10.715 -6.965 11.045 -6.635 ;
        RECT 9.355 -6.965 9.685 -6.635 ;
        RECT 7.995 -6.965 8.325 -6.635 ;
        RECT 6.635 -6.965 6.965 -6.635 ;
        RECT 5.275 -6.965 5.605 -6.635 ;
        RECT 3.915 -6.965 4.245 -6.635 ;
        RECT 2.555 -6.965 2.885 -6.635 ;
        RECT 1.195 -6.965 1.525 -6.635 ;
        RECT -0.165 -6.965 0.165 -6.635 ;
        RECT -1.525 -6.965 -1.195 -6.635 ;
        RECT 954.555 -6.965 954.885 -6.635 ;
        RECT 678.475 -6.96 954.885 -6.64 ;
        RECT 953.195 -6.965 953.525 -6.635 ;
        RECT 951.835 -6.965 952.165 -6.635 ;
        RECT 950.475 -6.965 950.805 -6.635 ;
        RECT 949.115 -6.965 949.445 -6.635 ;
        RECT 947.755 -6.965 948.085 -6.635 ;
        RECT 946.395 -6.965 946.725 -6.635 ;
        RECT 945.035 -6.965 945.365 -6.635 ;
        RECT 943.675 -6.965 944.005 -6.635 ;
        RECT 942.315 -6.965 942.645 -6.635 ;
        RECT 940.955 -6.965 941.285 -6.635 ;
        RECT 939.595 -6.965 939.925 -6.635 ;
        RECT 938.235 -6.965 938.565 -6.635 ;
        RECT 936.875 -6.965 937.205 -6.635 ;
        RECT 935.515 -6.965 935.845 -6.635 ;
        RECT 934.155 -6.965 934.485 -6.635 ;
        RECT 932.795 -6.965 933.125 -6.635 ;
        RECT 931.435 -6.965 931.765 -6.635 ;
        RECT 930.075 -6.965 930.405 -6.635 ;
        RECT 928.715 -6.965 929.045 -6.635 ;
        RECT 927.355 -6.965 927.685 -6.635 ;
        RECT 925.995 -6.965 926.325 -6.635 ;
        RECT 924.635 -6.965 924.965 -6.635 ;
        RECT 923.275 -6.965 923.605 -6.635 ;
        RECT 921.915 -6.965 922.245 -6.635 ;
        RECT 920.555 -6.965 920.885 -6.635 ;
        RECT 919.195 -6.965 919.525 -6.635 ;
        RECT 917.835 -6.965 918.165 -6.635 ;
        RECT 916.475 -6.965 916.805 -6.635 ;
        RECT 915.115 -6.965 915.445 -6.635 ;
        RECT 913.755 -6.965 914.085 -6.635 ;
        RECT 912.395 -6.965 912.725 -6.635 ;
        RECT 911.035 -6.965 911.365 -6.635 ;
        RECT 909.675 -6.965 910.005 -6.635 ;
        RECT 908.315 -6.965 908.645 -6.635 ;
        RECT 906.955 -6.965 907.285 -6.635 ;
        RECT 905.595 -6.965 905.925 -6.635 ;
        RECT 904.235 -6.965 904.565 -6.635 ;
        RECT 902.875 -6.965 903.205 -6.635 ;
        RECT 901.515 -6.965 901.845 -6.635 ;
        RECT 900.155 -6.965 900.485 -6.635 ;
        RECT 898.795 -6.965 899.125 -6.635 ;
        RECT 897.435 -6.965 897.765 -6.635 ;
        RECT 896.075 -6.965 896.405 -6.635 ;
        RECT 894.715 -6.965 895.045 -6.635 ;
        RECT 893.355 -6.965 893.685 -6.635 ;
        RECT 891.995 -6.965 892.325 -6.635 ;
        RECT 890.635 -6.965 890.965 -6.635 ;
        RECT 889.275 -6.965 889.605 -6.635 ;
        RECT 887.915 -6.965 888.245 -6.635 ;
        RECT 886.555 -6.965 886.885 -6.635 ;
        RECT 885.195 -6.965 885.525 -6.635 ;
        RECT 883.835 -6.965 884.165 -6.635 ;
        RECT 882.475 -6.965 882.805 -6.635 ;
        RECT 881.115 -6.965 881.445 -6.635 ;
        RECT 879.755 -6.965 880.085 -6.635 ;
        RECT 878.395 -6.965 878.725 -6.635 ;
        RECT 877.035 -6.965 877.365 -6.635 ;
        RECT 875.675 -6.965 876.005 -6.635 ;
        RECT 874.315 -6.965 874.645 -6.635 ;
        RECT 872.955 -6.965 873.285 -6.635 ;
        RECT 871.595 -6.965 871.925 -6.635 ;
        RECT 870.235 -6.965 870.565 -6.635 ;
        RECT 868.875 -6.965 869.205 -6.635 ;
        RECT 867.515 -6.965 867.845 -6.635 ;
        RECT 866.155 -6.965 866.485 -6.635 ;
        RECT 864.795 -6.965 865.125 -6.635 ;
        RECT 863.435 -6.965 863.765 -6.635 ;
        RECT 862.075 -6.965 862.405 -6.635 ;
        RECT 860.715 -6.965 861.045 -6.635 ;
        RECT 859.355 -6.965 859.685 -6.635 ;
        RECT 857.995 -6.965 858.325 -6.635 ;
        RECT 856.635 -6.965 856.965 -6.635 ;
        RECT 855.275 -6.965 855.605 -6.635 ;
        RECT 853.915 -6.965 854.245 -6.635 ;
        RECT 852.555 -6.965 852.885 -6.635 ;
        RECT 851.195 -6.965 851.525 -6.635 ;
        RECT 849.835 -6.965 850.165 -6.635 ;
        RECT 848.475 -6.965 848.805 -6.635 ;
        RECT 847.115 -6.965 847.445 -6.635 ;
        RECT 845.755 -6.965 846.085 -6.635 ;
        RECT 844.395 -6.965 844.725 -6.635 ;
        RECT 843.035 -6.965 843.365 -6.635 ;
        RECT 841.675 -6.965 842.005 -6.635 ;
        RECT 840.315 -6.965 840.645 -6.635 ;
        RECT 838.955 -6.965 839.285 -6.635 ;
        RECT 837.595 -6.965 837.925 -6.635 ;
        RECT 836.235 -6.965 836.565 -6.635 ;
        RECT 834.875 -6.965 835.205 -6.635 ;
        RECT 833.515 -6.965 833.845 -6.635 ;
        RECT 832.155 -6.965 832.485 -6.635 ;
        RECT 830.795 -6.965 831.125 -6.635 ;
        RECT 829.435 -6.965 829.765 -6.635 ;
        RECT 828.075 -6.965 828.405 -6.635 ;
        RECT 826.715 -6.965 827.045 -6.635 ;
        RECT 825.355 -6.965 825.685 -6.635 ;
        RECT 823.995 -6.965 824.325 -6.635 ;
        RECT 822.635 -6.965 822.965 -6.635 ;
        RECT 821.275 -6.965 821.605 -6.635 ;
        RECT 819.915 -6.965 820.245 -6.635 ;
        RECT 818.555 -6.965 818.885 -6.635 ;
        RECT 817.195 -6.965 817.525 -6.635 ;
        RECT 815.835 -6.965 816.165 -6.635 ;
        RECT 814.475 -6.965 814.805 -6.635 ;
        RECT 813.115 -6.965 813.445 -6.635 ;
        RECT 811.755 -6.965 812.085 -6.635 ;
        RECT 810.395 -6.965 810.725 -6.635 ;
        RECT 809.035 -6.965 809.365 -6.635 ;
        RECT 807.675 -6.965 808.005 -6.635 ;
        RECT 806.315 -6.965 806.645 -6.635 ;
        RECT 804.955 -6.965 805.285 -6.635 ;
        RECT 803.595 -6.965 803.925 -6.635 ;
        RECT 802.235 -6.965 802.565 -6.635 ;
        RECT 800.875 -6.965 801.205 -6.635 ;
        RECT 799.515 -6.965 799.845 -6.635 ;
        RECT 798.155 -6.965 798.485 -6.635 ;
        RECT 796.795 -6.965 797.125 -6.635 ;
        RECT 795.435 -6.965 795.765 -6.635 ;
        RECT 794.075 -6.965 794.405 -6.635 ;
        RECT 792.715 -6.965 793.045 -6.635 ;
        RECT 791.355 -6.965 791.685 -6.635 ;
        RECT 789.995 -6.965 790.325 -6.635 ;
        RECT 788.635 -6.965 788.965 -6.635 ;
        RECT 787.275 -6.965 787.605 -6.635 ;
        RECT 785.915 -6.965 786.245 -6.635 ;
        RECT 784.555 -6.965 784.885 -6.635 ;
        RECT 783.195 -6.965 783.525 -6.635 ;
        RECT 781.835 -6.965 782.165 -6.635 ;
        RECT 780.475 -6.965 780.805 -6.635 ;
        RECT 779.115 -6.965 779.445 -6.635 ;
        RECT 777.755 -6.965 778.085 -6.635 ;
        RECT 776.395 -6.965 776.725 -6.635 ;
        RECT 775.035 -6.965 775.365 -6.635 ;
        RECT 773.675 -6.965 774.005 -6.635 ;
        RECT 772.315 -6.965 772.645 -6.635 ;
        RECT 770.955 -6.965 771.285 -6.635 ;
        RECT 769.595 -6.965 769.925 -6.635 ;
        RECT 768.235 -6.965 768.565 -6.635 ;
        RECT 766.875 -6.965 767.205 -6.635 ;
        RECT 765.515 -6.965 765.845 -6.635 ;
        RECT 764.155 -6.965 764.485 -6.635 ;
        RECT 762.795 -6.965 763.125 -6.635 ;
        RECT 761.435 -6.965 761.765 -6.635 ;
        RECT 760.075 -6.965 760.405 -6.635 ;
        RECT 758.715 -6.965 759.045 -6.635 ;
        RECT 757.355 -6.965 757.685 -6.635 ;
        RECT 755.995 -6.965 756.325 -6.635 ;
        RECT 754.635 -6.965 754.965 -6.635 ;
        RECT 753.275 -6.965 753.605 -6.635 ;
        RECT 751.915 -6.965 752.245 -6.635 ;
        RECT 750.555 -6.965 750.885 -6.635 ;
        RECT 749.195 -6.965 749.525 -6.635 ;
        RECT 747.835 -6.965 748.165 -6.635 ;
        RECT 746.475 -6.965 746.805 -6.635 ;
        RECT 745.115 -6.965 745.445 -6.635 ;
        RECT 743.755 -6.965 744.085 -6.635 ;
        RECT 742.395 -6.965 742.725 -6.635 ;
        RECT 741.035 -6.965 741.365 -6.635 ;
        RECT 739.675 -6.965 740.005 -6.635 ;
        RECT 738.315 -6.965 738.645 -6.635 ;
        RECT 736.955 -6.965 737.285 -6.635 ;
        RECT 735.595 -6.965 735.925 -6.635 ;
        RECT 734.235 -6.965 734.565 -6.635 ;
        RECT 732.875 -6.965 733.205 -6.635 ;
        RECT 731.515 -6.965 731.845 -6.635 ;
        RECT 730.155 -6.965 730.485 -6.635 ;
        RECT 728.795 -6.965 729.125 -6.635 ;
        RECT 727.435 -6.965 727.765 -6.635 ;
        RECT 726.075 -6.965 726.405 -6.635 ;
        RECT 724.715 -6.965 725.045 -6.635 ;
        RECT 723.355 -6.965 723.685 -6.635 ;
        RECT 721.995 -6.965 722.325 -6.635 ;
        RECT 720.635 -6.965 720.965 -6.635 ;
        RECT 719.275 -6.965 719.605 -6.635 ;
        RECT 717.915 -6.965 718.245 -6.635 ;
        RECT 716.555 -6.965 716.885 -6.635 ;
        RECT 715.195 -6.965 715.525 -6.635 ;
        RECT 713.835 -6.965 714.165 -6.635 ;
        RECT 712.475 -6.965 712.805 -6.635 ;
        RECT 711.115 -6.965 711.445 -6.635 ;
        RECT 709.755 -6.965 710.085 -6.635 ;
        RECT 708.395 -6.965 708.725 -6.635 ;
        RECT 707.035 -6.965 707.365 -6.635 ;
        RECT 705.675 -6.965 706.005 -6.635 ;
        RECT 704.315 -6.965 704.645 -6.635 ;
        RECT 702.955 -6.965 703.285 -6.635 ;
        RECT 701.595 -6.965 701.925 -6.635 ;
        RECT 700.235 -6.965 700.565 -6.635 ;
        RECT 698.875 -6.965 699.205 -6.635 ;
        RECT 697.515 -6.965 697.845 -6.635 ;
        RECT 696.155 -6.965 696.485 -6.635 ;
        RECT 694.795 -6.965 695.125 -6.635 ;
        RECT 693.435 -6.965 693.765 -6.635 ;
        RECT 692.075 -6.965 692.405 -6.635 ;
        RECT 690.715 -6.965 691.045 -6.635 ;
        RECT 689.355 -6.965 689.685 -6.635 ;
        RECT 687.995 -6.965 688.325 -6.635 ;
        RECT 686.635 -6.965 686.965 -6.635 ;
        RECT 685.275 -6.965 685.605 -6.635 ;
        RECT 683.915 -6.965 684.245 -6.635 ;
        RECT 682.555 -6.965 682.885 -6.635 ;
        RECT 681.195 -6.965 681.525 -6.635 ;
        RECT 679.835 -6.965 680.165 -6.635 ;
        RECT 678.475 -6.965 678.805 -6.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.275 -8.325 651.605 -7.995 ;
        RECT 649.915 -8.325 650.245 -7.995 ;
        RECT 648.555 -8.325 648.885 -7.995 ;
        RECT 647.195 -8.325 647.525 -7.995 ;
        RECT 645.835 -8.325 646.165 -7.995 ;
        RECT 644.475 -8.325 644.805 -7.995 ;
        RECT 643.115 -8.325 643.445 -7.995 ;
        RECT 641.755 -8.325 642.085 -7.995 ;
        RECT 640.395 -8.325 640.725 -7.995 ;
        RECT 639.035 -8.325 639.365 -7.995 ;
        RECT 637.675 -8.325 638.005 -7.995 ;
        RECT 636.315 -8.325 636.645 -7.995 ;
        RECT 634.955 -8.325 635.285 -7.995 ;
        RECT 633.595 -8.325 633.925 -7.995 ;
        RECT 632.235 -8.325 632.565 -7.995 ;
        RECT 630.875 -8.325 631.205 -7.995 ;
        RECT 629.515 -8.325 629.845 -7.995 ;
        RECT 628.155 -8.325 628.485 -7.995 ;
        RECT 626.795 -8.325 627.125 -7.995 ;
        RECT 625.435 -8.325 625.765 -7.995 ;
        RECT 624.075 -8.325 624.405 -7.995 ;
        RECT 622.715 -8.325 623.045 -7.995 ;
        RECT 621.355 -8.325 621.685 -7.995 ;
        RECT 619.995 -8.325 620.325 -7.995 ;
        RECT 618.635 -8.325 618.965 -7.995 ;
        RECT 617.275 -8.325 617.605 -7.995 ;
        RECT 615.915 -8.325 616.245 -7.995 ;
        RECT 614.555 -8.325 614.885 -7.995 ;
        RECT 613.195 -8.325 613.525 -7.995 ;
        RECT 611.835 -8.325 612.165 -7.995 ;
        RECT 610.475 -8.325 610.805 -7.995 ;
        RECT 609.115 -8.325 609.445 -7.995 ;
        RECT 607.755 -8.325 608.085 -7.995 ;
        RECT 606.395 -8.325 606.725 -7.995 ;
        RECT 605.035 -8.325 605.365 -7.995 ;
        RECT 603.675 -8.325 604.005 -7.995 ;
        RECT 602.315 -8.325 602.645 -7.995 ;
        RECT 600.955 -8.325 601.285 -7.995 ;
        RECT 599.595 -8.325 599.925 -7.995 ;
        RECT 598.235 -8.325 598.565 -7.995 ;
        RECT 596.875 -8.325 597.205 -7.995 ;
        RECT 595.515 -8.325 595.845 -7.995 ;
        RECT 594.155 -8.325 594.485 -7.995 ;
        RECT 592.795 -8.325 593.125 -7.995 ;
        RECT 591.435 -8.325 591.765 -7.995 ;
        RECT 590.075 -8.325 590.405 -7.995 ;
        RECT 588.715 -8.325 589.045 -7.995 ;
        RECT 587.355 -8.325 587.685 -7.995 ;
        RECT 585.995 -8.325 586.325 -7.995 ;
        RECT 584.635 -8.325 584.965 -7.995 ;
        RECT 583.275 -8.325 583.605 -7.995 ;
        RECT 581.915 -8.325 582.245 -7.995 ;
        RECT 580.555 -8.325 580.885 -7.995 ;
        RECT 579.195 -8.325 579.525 -7.995 ;
        RECT 577.835 -8.325 578.165 -7.995 ;
        RECT 576.475 -8.325 576.805 -7.995 ;
        RECT 575.115 -8.325 575.445 -7.995 ;
        RECT 573.755 -8.325 574.085 -7.995 ;
        RECT 572.395 -8.325 572.725 -7.995 ;
        RECT 571.035 -8.325 571.365 -7.995 ;
        RECT 569.675 -8.325 570.005 -7.995 ;
        RECT 568.315 -8.325 568.645 -7.995 ;
        RECT 566.955 -8.325 567.285 -7.995 ;
        RECT 565.595 -8.325 565.925 -7.995 ;
        RECT 564.235 -8.325 564.565 -7.995 ;
        RECT 562.875 -8.325 563.205 -7.995 ;
        RECT 561.515 -8.325 561.845 -7.995 ;
        RECT 560.155 -8.325 560.485 -7.995 ;
        RECT 558.795 -8.325 559.125 -7.995 ;
        RECT 557.435 -8.325 557.765 -7.995 ;
        RECT 556.075 -8.325 556.405 -7.995 ;
        RECT 554.715 -8.325 555.045 -7.995 ;
        RECT 553.355 -8.325 553.685 -7.995 ;
        RECT 551.995 -8.325 552.325 -7.995 ;
        RECT 550.635 -8.325 550.965 -7.995 ;
        RECT 549.275 -8.325 549.605 -7.995 ;
        RECT 547.915 -8.325 548.245 -7.995 ;
        RECT 546.555 -8.325 546.885 -7.995 ;
        RECT 545.195 -8.325 545.525 -7.995 ;
        RECT 543.835 -8.325 544.165 -7.995 ;
        RECT 542.475 -8.325 542.805 -7.995 ;
        RECT 541.115 -8.325 541.445 -7.995 ;
        RECT 539.755 -8.325 540.085 -7.995 ;
        RECT 538.395 -8.325 538.725 -7.995 ;
        RECT 537.035 -8.325 537.365 -7.995 ;
        RECT 535.675 -8.325 536.005 -7.995 ;
        RECT 534.315 -8.325 534.645 -7.995 ;
        RECT 532.955 -8.325 533.285 -7.995 ;
        RECT 531.595 -8.325 531.925 -7.995 ;
        RECT 530.235 -8.325 530.565 -7.995 ;
        RECT 528.875 -8.325 529.205 -7.995 ;
        RECT 527.515 -8.325 527.845 -7.995 ;
        RECT 526.155 -8.325 526.485 -7.995 ;
        RECT 524.795 -8.325 525.125 -7.995 ;
        RECT 523.435 -8.325 523.765 -7.995 ;
        RECT 522.075 -8.325 522.405 -7.995 ;
        RECT 520.715 -8.325 521.045 -7.995 ;
        RECT 519.355 -8.325 519.685 -7.995 ;
        RECT 517.995 -8.325 518.325 -7.995 ;
        RECT 516.635 -8.325 516.965 -7.995 ;
        RECT 515.275 -8.325 515.605 -7.995 ;
        RECT 513.915 -8.325 514.245 -7.995 ;
        RECT 512.555 -8.325 512.885 -7.995 ;
        RECT 511.195 -8.325 511.525 -7.995 ;
        RECT 509.835 -8.325 510.165 -7.995 ;
        RECT 508.475 -8.325 508.805 -7.995 ;
        RECT 507.115 -8.325 507.445 -7.995 ;
        RECT 505.755 -8.325 506.085 -7.995 ;
        RECT 504.395 -8.325 504.725 -7.995 ;
        RECT 503.035 -8.325 503.365 -7.995 ;
        RECT 501.675 -8.325 502.005 -7.995 ;
        RECT 500.315 -8.325 500.645 -7.995 ;
        RECT 498.955 -8.325 499.285 -7.995 ;
        RECT 497.595 -8.325 497.925 -7.995 ;
        RECT 496.235 -8.325 496.565 -7.995 ;
        RECT 494.875 -8.325 495.205 -7.995 ;
        RECT 493.515 -8.325 493.845 -7.995 ;
        RECT 492.155 -8.325 492.485 -7.995 ;
        RECT 490.795 -8.325 491.125 -7.995 ;
        RECT 489.435 -8.325 489.765 -7.995 ;
        RECT 488.075 -8.325 488.405 -7.995 ;
        RECT 486.715 -8.325 487.045 -7.995 ;
        RECT 485.355 -8.325 485.685 -7.995 ;
        RECT 483.995 -8.325 484.325 -7.995 ;
        RECT 482.635 -8.325 482.965 -7.995 ;
        RECT 481.275 -8.325 481.605 -7.995 ;
        RECT 479.915 -8.325 480.245 -7.995 ;
        RECT 478.555 -8.325 478.885 -7.995 ;
        RECT 477.195 -8.325 477.525 -7.995 ;
        RECT 475.835 -8.325 476.165 -7.995 ;
        RECT 474.475 -8.325 474.805 -7.995 ;
        RECT 473.115 -8.325 473.445 -7.995 ;
        RECT 471.755 -8.325 472.085 -7.995 ;
        RECT 470.395 -8.325 470.725 -7.995 ;
        RECT 469.035 -8.325 469.365 -7.995 ;
        RECT 467.675 -8.325 468.005 -7.995 ;
        RECT 466.315 -8.325 466.645 -7.995 ;
        RECT 464.955 -8.325 465.285 -7.995 ;
        RECT 463.595 -8.325 463.925 -7.995 ;
        RECT 462.235 -8.325 462.565 -7.995 ;
        RECT 460.875 -8.325 461.205 -7.995 ;
        RECT 459.515 -8.325 459.845 -7.995 ;
        RECT 458.155 -8.325 458.485 -7.995 ;
        RECT 456.795 -8.325 457.125 -7.995 ;
        RECT 455.435 -8.325 455.765 -7.995 ;
        RECT 454.075 -8.325 454.405 -7.995 ;
        RECT 452.715 -8.325 453.045 -7.995 ;
        RECT 451.355 -8.325 451.685 -7.995 ;
        RECT 449.995 -8.325 450.325 -7.995 ;
        RECT 448.635 -8.325 448.965 -7.995 ;
        RECT 447.275 -8.325 447.605 -7.995 ;
        RECT 445.915 -8.325 446.245 -7.995 ;
        RECT 444.555 -8.325 444.885 -7.995 ;
        RECT 443.195 -8.325 443.525 -7.995 ;
        RECT 441.835 -8.325 442.165 -7.995 ;
        RECT 440.475 -8.325 440.805 -7.995 ;
        RECT 439.115 -8.325 439.445 -7.995 ;
        RECT 437.755 -8.325 438.085 -7.995 ;
        RECT 436.395 -8.325 436.725 -7.995 ;
        RECT 435.035 -8.325 435.365 -7.995 ;
        RECT 433.675 -8.325 434.005 -7.995 ;
        RECT 432.315 -8.325 432.645 -7.995 ;
        RECT 430.955 -8.325 431.285 -7.995 ;
        RECT 429.595 -8.325 429.925 -7.995 ;
        RECT 428.235 -8.325 428.565 -7.995 ;
        RECT 426.875 -8.325 427.205 -7.995 ;
        RECT 425.515 -8.325 425.845 -7.995 ;
        RECT 424.155 -8.325 424.485 -7.995 ;
        RECT 422.795 -8.325 423.125 -7.995 ;
        RECT 421.435 -8.325 421.765 -7.995 ;
        RECT 420.075 -8.325 420.405 -7.995 ;
        RECT 418.715 -8.325 419.045 -7.995 ;
        RECT 417.355 -8.325 417.685 -7.995 ;
        RECT 415.995 -8.325 416.325 -7.995 ;
        RECT 414.635 -8.325 414.965 -7.995 ;
        RECT 413.275 -8.325 413.605 -7.995 ;
        RECT 411.915 -8.325 412.245 -7.995 ;
        RECT 410.555 -8.325 410.885 -7.995 ;
        RECT 409.195 -8.325 409.525 -7.995 ;
        RECT 407.835 -8.325 408.165 -7.995 ;
        RECT 406.475 -8.325 406.805 -7.995 ;
        RECT 405.115 -8.325 405.445 -7.995 ;
        RECT 403.755 -8.325 404.085 -7.995 ;
        RECT 402.395 -8.325 402.725 -7.995 ;
        RECT 401.035 -8.325 401.365 -7.995 ;
        RECT 399.675 -8.325 400.005 -7.995 ;
        RECT 398.315 -8.325 398.645 -7.995 ;
        RECT 396.955 -8.325 397.285 -7.995 ;
        RECT 395.595 -8.325 395.925 -7.995 ;
        RECT 394.235 -8.325 394.565 -7.995 ;
        RECT 392.875 -8.325 393.205 -7.995 ;
        RECT 391.515 -8.325 391.845 -7.995 ;
        RECT 390.155 -8.325 390.485 -7.995 ;
        RECT 388.795 -8.325 389.125 -7.995 ;
        RECT 387.435 -8.325 387.765 -7.995 ;
        RECT 386.075 -8.325 386.405 -7.995 ;
        RECT 384.715 -8.325 385.045 -7.995 ;
        RECT 383.355 -8.325 383.685 -7.995 ;
        RECT 381.995 -8.325 382.325 -7.995 ;
        RECT 380.635 -8.325 380.965 -7.995 ;
        RECT 379.275 -8.325 379.605 -7.995 ;
        RECT 377.915 -8.325 378.245 -7.995 ;
        RECT 376.555 -8.325 376.885 -7.995 ;
        RECT 375.195 -8.325 375.525 -7.995 ;
        RECT 373.835 -8.325 374.165 -7.995 ;
        RECT 372.475 -8.325 372.805 -7.995 ;
        RECT 371.115 -8.325 371.445 -7.995 ;
        RECT 369.755 -8.325 370.085 -7.995 ;
        RECT 368.395 -8.325 368.725 -7.995 ;
        RECT 367.035 -8.325 367.365 -7.995 ;
        RECT 365.675 -8.325 366.005 -7.995 ;
        RECT 364.315 -8.325 364.645 -7.995 ;
        RECT 362.955 -8.325 363.285 -7.995 ;
        RECT 361.595 -8.325 361.925 -7.995 ;
        RECT 360.235 -8.325 360.565 -7.995 ;
        RECT 358.875 -8.325 359.205 -7.995 ;
        RECT 357.515 -8.325 357.845 -7.995 ;
        RECT 356.155 -8.325 356.485 -7.995 ;
        RECT 354.795 -8.325 355.125 -7.995 ;
        RECT 353.435 -8.325 353.765 -7.995 ;
        RECT 352.075 -8.325 352.405 -7.995 ;
        RECT 350.715 -8.325 351.045 -7.995 ;
        RECT 349.355 -8.325 349.685 -7.995 ;
        RECT 347.995 -8.325 348.325 -7.995 ;
        RECT 346.635 -8.325 346.965 -7.995 ;
        RECT 345.275 -8.325 345.605 -7.995 ;
        RECT 343.915 -8.325 344.245 -7.995 ;
        RECT 342.555 -8.325 342.885 -7.995 ;
        RECT 341.195 -8.325 341.525 -7.995 ;
        RECT 339.835 -8.325 340.165 -7.995 ;
        RECT 338.475 -8.325 338.805 -7.995 ;
        RECT 337.115 -8.325 337.445 -7.995 ;
        RECT 335.755 -8.325 336.085 -7.995 ;
        RECT 334.395 -8.325 334.725 -7.995 ;
        RECT 333.035 -8.325 333.365 -7.995 ;
        RECT 331.675 -8.325 332.005 -7.995 ;
        RECT 330.315 -8.325 330.645 -7.995 ;
        RECT 328.955 -8.325 329.285 -7.995 ;
        RECT 327.595 -8.325 327.925 -7.995 ;
        RECT 326.235 -8.325 326.565 -7.995 ;
        RECT 324.875 -8.325 325.205 -7.995 ;
        RECT 323.515 -8.325 323.845 -7.995 ;
        RECT 322.155 -8.325 322.485 -7.995 ;
        RECT 320.795 -8.325 321.125 -7.995 ;
        RECT 319.435 -8.325 319.765 -7.995 ;
        RECT 318.075 -8.325 318.405 -7.995 ;
        RECT 316.715 -8.325 317.045 -7.995 ;
        RECT 315.355 -8.325 315.685 -7.995 ;
        RECT 313.995 -8.325 314.325 -7.995 ;
        RECT 312.635 -8.325 312.965 -7.995 ;
        RECT 311.275 -8.325 311.605 -7.995 ;
        RECT 309.915 -8.325 310.245 -7.995 ;
        RECT 308.555 -8.325 308.885 -7.995 ;
        RECT 307.195 -8.325 307.525 -7.995 ;
        RECT 305.835 -8.325 306.165 -7.995 ;
        RECT 304.475 -8.325 304.805 -7.995 ;
        RECT 303.115 -8.325 303.445 -7.995 ;
        RECT 301.755 -8.325 302.085 -7.995 ;
        RECT 300.395 -8.325 300.725 -7.995 ;
        RECT 299.035 -8.325 299.365 -7.995 ;
        RECT 297.675 -8.325 298.005 -7.995 ;
        RECT 296.315 -8.325 296.645 -7.995 ;
        RECT 294.955 -8.325 295.285 -7.995 ;
        RECT 293.595 -8.325 293.925 -7.995 ;
        RECT 292.235 -8.325 292.565 -7.995 ;
        RECT 290.875 -8.325 291.205 -7.995 ;
        RECT 289.515 -8.325 289.845 -7.995 ;
        RECT 288.155 -8.325 288.485 -7.995 ;
        RECT 286.795 -8.325 287.125 -7.995 ;
        RECT 285.435 -8.325 285.765 -7.995 ;
        RECT 284.075 -8.325 284.405 -7.995 ;
        RECT 282.715 -8.325 283.045 -7.995 ;
        RECT 281.355 -8.325 281.685 -7.995 ;
        RECT 279.995 -8.325 280.325 -7.995 ;
        RECT 278.635 -8.325 278.965 -7.995 ;
        RECT 277.275 -8.325 277.605 -7.995 ;
        RECT 275.915 -8.325 276.245 -7.995 ;
        RECT 274.555 -8.325 274.885 -7.995 ;
        RECT 273.195 -8.325 273.525 -7.995 ;
        RECT 271.835 -8.325 272.165 -7.995 ;
        RECT 270.475 -8.325 270.805 -7.995 ;
        RECT 269.115 -8.325 269.445 -7.995 ;
        RECT 267.755 -8.325 268.085 -7.995 ;
        RECT 266.395 -8.325 266.725 -7.995 ;
        RECT 265.035 -8.325 265.365 -7.995 ;
        RECT 263.675 -8.325 264.005 -7.995 ;
        RECT 262.315 -8.325 262.645 -7.995 ;
        RECT 260.955 -8.325 261.285 -7.995 ;
        RECT 259.595 -8.325 259.925 -7.995 ;
        RECT 258.235 -8.325 258.565 -7.995 ;
        RECT 256.875 -8.325 257.205 -7.995 ;
        RECT 255.515 -8.325 255.845 -7.995 ;
        RECT 254.155 -8.325 254.485 -7.995 ;
        RECT 252.795 -8.325 253.125 -7.995 ;
        RECT 251.435 -8.325 251.765 -7.995 ;
        RECT 250.075 -8.325 250.405 -7.995 ;
        RECT 248.715 -8.325 249.045 -7.995 ;
        RECT 247.355 -8.325 247.685 -7.995 ;
        RECT 245.995 -8.325 246.325 -7.995 ;
        RECT 244.635 -8.325 244.965 -7.995 ;
        RECT 243.275 -8.325 243.605 -7.995 ;
        RECT 241.915 -8.325 242.245 -7.995 ;
        RECT 240.555 -8.325 240.885 -7.995 ;
        RECT 239.195 -8.325 239.525 -7.995 ;
        RECT 237.835 -8.325 238.165 -7.995 ;
        RECT 236.475 -8.325 236.805 -7.995 ;
        RECT 235.115 -8.325 235.445 -7.995 ;
        RECT 233.755 -8.325 234.085 -7.995 ;
        RECT 232.395 -8.325 232.725 -7.995 ;
        RECT 231.035 -8.325 231.365 -7.995 ;
        RECT 229.675 -8.325 230.005 -7.995 ;
        RECT 228.315 -8.325 228.645 -7.995 ;
        RECT 226.955 -8.325 227.285 -7.995 ;
        RECT 225.595 -8.325 225.925 -7.995 ;
        RECT 224.235 -8.325 224.565 -7.995 ;
        RECT 222.875 -8.325 223.205 -7.995 ;
        RECT 221.515 -8.325 221.845 -7.995 ;
        RECT 220.155 -8.325 220.485 -7.995 ;
        RECT 218.795 -8.325 219.125 -7.995 ;
        RECT 217.435 -8.325 217.765 -7.995 ;
        RECT 216.075 -8.325 216.405 -7.995 ;
        RECT 214.715 -8.325 215.045 -7.995 ;
        RECT 213.355 -8.325 213.685 -7.995 ;
        RECT 211.995 -8.325 212.325 -7.995 ;
        RECT 210.635 -8.325 210.965 -7.995 ;
        RECT 209.275 -8.325 209.605 -7.995 ;
        RECT 207.915 -8.325 208.245 -7.995 ;
        RECT 206.555 -8.325 206.885 -7.995 ;
        RECT 205.195 -8.325 205.525 -7.995 ;
        RECT 203.835 -8.325 204.165 -7.995 ;
        RECT 202.475 -8.325 202.805 -7.995 ;
        RECT 201.115 -8.325 201.445 -7.995 ;
        RECT 199.755 -8.325 200.085 -7.995 ;
        RECT 198.395 -8.325 198.725 -7.995 ;
        RECT 197.035 -8.325 197.365 -7.995 ;
        RECT 195.675 -8.325 196.005 -7.995 ;
        RECT 194.315 -8.325 194.645 -7.995 ;
        RECT 192.955 -8.325 193.285 -7.995 ;
        RECT 191.595 -8.325 191.925 -7.995 ;
        RECT 190.235 -8.325 190.565 -7.995 ;
        RECT 188.875 -8.325 189.205 -7.995 ;
        RECT 187.515 -8.325 187.845 -7.995 ;
        RECT 186.155 -8.325 186.485 -7.995 ;
        RECT 184.795 -8.325 185.125 -7.995 ;
        RECT 183.435 -8.325 183.765 -7.995 ;
        RECT 182.075 -8.325 182.405 -7.995 ;
        RECT 180.715 -8.325 181.045 -7.995 ;
        RECT 179.355 -8.325 179.685 -7.995 ;
        RECT 177.995 -8.325 178.325 -7.995 ;
        RECT 176.635 -8.325 176.965 -7.995 ;
        RECT 175.275 -8.325 175.605 -7.995 ;
        RECT 173.915 -8.325 174.245 -7.995 ;
        RECT 172.555 -8.325 172.885 -7.995 ;
        RECT 171.195 -8.325 171.525 -7.995 ;
        RECT 169.835 -8.325 170.165 -7.995 ;
        RECT 168.475 -8.325 168.805 -7.995 ;
        RECT 167.115 -8.325 167.445 -7.995 ;
        RECT 165.755 -8.325 166.085 -7.995 ;
        RECT 164.395 -8.325 164.725 -7.995 ;
        RECT 163.035 -8.325 163.365 -7.995 ;
        RECT 161.675 -8.325 162.005 -7.995 ;
        RECT 160.315 -8.325 160.645 -7.995 ;
        RECT 158.955 -8.325 159.285 -7.995 ;
        RECT 157.595 -8.325 157.925 -7.995 ;
        RECT 156.235 -8.325 156.565 -7.995 ;
        RECT 154.875 -8.325 155.205 -7.995 ;
        RECT 153.515 -8.325 153.845 -7.995 ;
        RECT 152.155 -8.325 152.485 -7.995 ;
        RECT 150.795 -8.325 151.125 -7.995 ;
        RECT 149.435 -8.325 149.765 -7.995 ;
        RECT 148.075 -8.325 148.405 -7.995 ;
        RECT 146.715 -8.325 147.045 -7.995 ;
        RECT 145.355 -8.325 145.685 -7.995 ;
        RECT 143.995 -8.325 144.325 -7.995 ;
        RECT 142.635 -8.325 142.965 -7.995 ;
        RECT 141.275 -8.325 141.605 -7.995 ;
        RECT 139.915 -8.325 140.245 -7.995 ;
        RECT 138.555 -8.325 138.885 -7.995 ;
        RECT 137.195 -8.325 137.525 -7.995 ;
        RECT 135.835 -8.325 136.165 -7.995 ;
        RECT 134.475 -8.325 134.805 -7.995 ;
        RECT 133.115 -8.325 133.445 -7.995 ;
        RECT 131.755 -8.325 132.085 -7.995 ;
        RECT 130.395 -8.325 130.725 -7.995 ;
        RECT 129.035 -8.325 129.365 -7.995 ;
        RECT 127.675 -8.325 128.005 -7.995 ;
        RECT 126.315 -8.325 126.645 -7.995 ;
        RECT 124.955 -8.325 125.285 -7.995 ;
        RECT 123.595 -8.325 123.925 -7.995 ;
        RECT 122.235 -8.325 122.565 -7.995 ;
        RECT 120.875 -8.325 121.205 -7.995 ;
        RECT 119.515 -8.325 119.845 -7.995 ;
        RECT 118.155 -8.325 118.485 -7.995 ;
        RECT 116.795 -8.325 117.125 -7.995 ;
        RECT 115.435 -8.325 115.765 -7.995 ;
        RECT 114.075 -8.325 114.405 -7.995 ;
        RECT 112.715 -8.325 113.045 -7.995 ;
        RECT 111.355 -8.325 111.685 -7.995 ;
        RECT 109.995 -8.325 110.325 -7.995 ;
        RECT 108.635 -8.325 108.965 -7.995 ;
        RECT 107.275 -8.325 107.605 -7.995 ;
        RECT 105.915 -8.325 106.245 -7.995 ;
        RECT 104.555 -8.325 104.885 -7.995 ;
        RECT 103.195 -8.325 103.525 -7.995 ;
        RECT 101.835 -8.325 102.165 -7.995 ;
        RECT 100.475 -8.325 100.805 -7.995 ;
        RECT 99.115 -8.325 99.445 -7.995 ;
        RECT 97.755 -8.325 98.085 -7.995 ;
        RECT 96.395 -8.325 96.725 -7.995 ;
        RECT 95.035 -8.325 95.365 -7.995 ;
        RECT 93.675 -8.325 94.005 -7.995 ;
        RECT 92.315 -8.325 92.645 -7.995 ;
        RECT 90.955 -8.325 91.285 -7.995 ;
        RECT 89.595 -8.325 89.925 -7.995 ;
        RECT 88.235 -8.325 88.565 -7.995 ;
        RECT 86.875 -8.325 87.205 -7.995 ;
        RECT 85.515 -8.325 85.845 -7.995 ;
        RECT 84.155 -8.325 84.485 -7.995 ;
        RECT 82.795 -8.325 83.125 -7.995 ;
        RECT 81.435 -8.325 81.765 -7.995 ;
        RECT 80.075 -8.325 80.405 -7.995 ;
        RECT 78.715 -8.325 79.045 -7.995 ;
        RECT 77.355 -8.325 77.685 -7.995 ;
        RECT 75.995 -8.325 76.325 -7.995 ;
        RECT 74.635 -8.325 74.965 -7.995 ;
        RECT 73.275 -8.325 73.605 -7.995 ;
        RECT 71.915 -8.325 72.245 -7.995 ;
        RECT 70.555 -8.325 70.885 -7.995 ;
        RECT 69.195 -8.325 69.525 -7.995 ;
        RECT 67.835 -8.325 68.165 -7.995 ;
        RECT 66.475 -8.325 66.805 -7.995 ;
        RECT 65.115 -8.325 65.445 -7.995 ;
        RECT 63.755 -8.325 64.085 -7.995 ;
        RECT 62.395 -8.325 62.725 -7.995 ;
        RECT 61.035 -8.325 61.365 -7.995 ;
        RECT 59.675 -8.325 60.005 -7.995 ;
        RECT 58.315 -8.325 58.645 -7.995 ;
        RECT 56.955 -8.325 57.285 -7.995 ;
        RECT 55.595 -8.325 55.925 -7.995 ;
        RECT 54.235 -8.325 54.565 -7.995 ;
        RECT 52.875 -8.325 53.205 -7.995 ;
        RECT 51.515 -8.325 51.845 -7.995 ;
        RECT 50.155 -8.325 50.485 -7.995 ;
        RECT 48.795 -8.325 49.125 -7.995 ;
        RECT 47.435 -8.325 47.765 -7.995 ;
        RECT 46.075 -8.325 46.405 -7.995 ;
        RECT 44.715 -8.325 45.045 -7.995 ;
        RECT 43.355 -8.325 43.685 -7.995 ;
        RECT 41.995 -8.325 42.325 -7.995 ;
        RECT 40.635 -8.325 40.965 -7.995 ;
        RECT 39.275 -8.325 39.605 -7.995 ;
        RECT 37.915 -8.325 38.245 -7.995 ;
        RECT 36.555 -8.325 36.885 -7.995 ;
        RECT 35.195 -8.325 35.525 -7.995 ;
        RECT 33.835 -8.325 34.165 -7.995 ;
        RECT 32.475 -8.325 32.805 -7.995 ;
        RECT 31.115 -8.325 31.445 -7.995 ;
        RECT 29.755 -8.325 30.085 -7.995 ;
        RECT 28.395 -8.325 28.725 -7.995 ;
        RECT 27.035 -8.325 27.365 -7.995 ;
        RECT 25.675 -8.325 26.005 -7.995 ;
        RECT 24.315 -8.325 24.645 -7.995 ;
        RECT 22.955 -8.325 23.285 -7.995 ;
        RECT 21.595 -8.325 21.925 -7.995 ;
        RECT 20.235 -8.325 20.565 -7.995 ;
        RECT 18.875 -8.325 19.205 -7.995 ;
        RECT 17.515 -8.325 17.845 -7.995 ;
        RECT 16.155 -8.325 16.485 -7.995 ;
        RECT 14.795 -8.325 15.125 -7.995 ;
        RECT 13.435 -8.325 13.765 -7.995 ;
        RECT 12.075 -8.325 12.405 -7.995 ;
        RECT 10.715 -8.325 11.045 -7.995 ;
        RECT 9.355 -8.325 9.685 -7.995 ;
        RECT 7.995 -8.325 8.325 -7.995 ;
        RECT 6.635 -8.325 6.965 -7.995 ;
        RECT 5.275 -8.325 5.605 -7.995 ;
        RECT 3.915 -8.325 4.245 -7.995 ;
        RECT 2.555 -8.325 2.885 -7.995 ;
        RECT 1.195 -8.325 1.525 -7.995 ;
        RECT -0.165 -8.325 0.165 -7.995 ;
        RECT -1.525 -8.325 -1.195 -7.995 ;
        RECT -1.525 -8.32 678.475 -8 ;
        RECT 677.115 -8.325 677.445 -7.995 ;
        RECT 675.755 -8.325 676.085 -7.995 ;
        RECT 674.395 -8.325 674.725 -7.995 ;
        RECT 673.035 -8.325 673.365 -7.995 ;
        RECT 671.675 -8.325 672.005 -7.995 ;
        RECT 670.315 -8.325 670.645 -7.995 ;
        RECT 668.955 -8.325 669.285 -7.995 ;
        RECT 667.595 -8.325 667.925 -7.995 ;
        RECT 666.235 -8.325 666.565 -7.995 ;
        RECT 664.875 -8.325 665.205 -7.995 ;
        RECT 663.515 -8.325 663.845 -7.995 ;
        RECT 662.155 -8.325 662.485 -7.995 ;
        RECT 660.795 -8.325 661.125 -7.995 ;
        RECT 659.435 -8.325 659.765 -7.995 ;
        RECT 658.075 -8.325 658.405 -7.995 ;
        RECT 656.715 -8.325 657.045 -7.995 ;
        RECT 655.355 -8.325 655.685 -7.995 ;
        RECT 653.995 -8.325 654.325 -7.995 ;
        RECT 652.635 -8.325 652.965 -7.995 ;
        RECT 954.555 -8.325 954.885 -7.995 ;
        RECT 678.475 -8.32 954.885 -8 ;
        RECT 953.195 -8.325 953.525 -7.995 ;
        RECT 951.835 -8.325 952.165 -7.995 ;
        RECT 950.475 -8.325 950.805 -7.995 ;
        RECT 949.115 -8.325 949.445 -7.995 ;
        RECT 947.755 -8.325 948.085 -7.995 ;
        RECT 946.395 -8.325 946.725 -7.995 ;
        RECT 945.035 -8.325 945.365 -7.995 ;
        RECT 943.675 -8.325 944.005 -7.995 ;
        RECT 942.315 -8.325 942.645 -7.995 ;
        RECT 940.955 -8.325 941.285 -7.995 ;
        RECT 939.595 -8.325 939.925 -7.995 ;
        RECT 938.235 -8.325 938.565 -7.995 ;
        RECT 936.875 -8.325 937.205 -7.995 ;
        RECT 935.515 -8.325 935.845 -7.995 ;
        RECT 934.155 -8.325 934.485 -7.995 ;
        RECT 932.795 -8.325 933.125 -7.995 ;
        RECT 931.435 -8.325 931.765 -7.995 ;
        RECT 930.075 -8.325 930.405 -7.995 ;
        RECT 928.715 -8.325 929.045 -7.995 ;
        RECT 927.355 -8.325 927.685 -7.995 ;
        RECT 925.995 -8.325 926.325 -7.995 ;
        RECT 924.635 -8.325 924.965 -7.995 ;
        RECT 923.275 -8.325 923.605 -7.995 ;
        RECT 921.915 -8.325 922.245 -7.995 ;
        RECT 920.555 -8.325 920.885 -7.995 ;
        RECT 919.195 -8.325 919.525 -7.995 ;
        RECT 917.835 -8.325 918.165 -7.995 ;
        RECT 916.475 -8.325 916.805 -7.995 ;
        RECT 915.115 -8.325 915.445 -7.995 ;
        RECT 913.755 -8.325 914.085 -7.995 ;
        RECT 912.395 -8.325 912.725 -7.995 ;
        RECT 911.035 -8.325 911.365 -7.995 ;
        RECT 909.675 -8.325 910.005 -7.995 ;
        RECT 908.315 -8.325 908.645 -7.995 ;
        RECT 906.955 -8.325 907.285 -7.995 ;
        RECT 905.595 -8.325 905.925 -7.995 ;
        RECT 904.235 -8.325 904.565 -7.995 ;
        RECT 902.875 -8.325 903.205 -7.995 ;
        RECT 901.515 -8.325 901.845 -7.995 ;
        RECT 900.155 -8.325 900.485 -7.995 ;
        RECT 898.795 -8.325 899.125 -7.995 ;
        RECT 897.435 -8.325 897.765 -7.995 ;
        RECT 896.075 -8.325 896.405 -7.995 ;
        RECT 894.715 -8.325 895.045 -7.995 ;
        RECT 893.355 -8.325 893.685 -7.995 ;
        RECT 891.995 -8.325 892.325 -7.995 ;
        RECT 890.635 -8.325 890.965 -7.995 ;
        RECT 889.275 -8.325 889.605 -7.995 ;
        RECT 887.915 -8.325 888.245 -7.995 ;
        RECT 886.555 -8.325 886.885 -7.995 ;
        RECT 885.195 -8.325 885.525 -7.995 ;
        RECT 883.835 -8.325 884.165 -7.995 ;
        RECT 882.475 -8.325 882.805 -7.995 ;
        RECT 881.115 -8.325 881.445 -7.995 ;
        RECT 879.755 -8.325 880.085 -7.995 ;
        RECT 878.395 -8.325 878.725 -7.995 ;
        RECT 877.035 -8.325 877.365 -7.995 ;
        RECT 875.675 -8.325 876.005 -7.995 ;
        RECT 874.315 -8.325 874.645 -7.995 ;
        RECT 872.955 -8.325 873.285 -7.995 ;
        RECT 871.595 -8.325 871.925 -7.995 ;
        RECT 870.235 -8.325 870.565 -7.995 ;
        RECT 868.875 -8.325 869.205 -7.995 ;
        RECT 867.515 -8.325 867.845 -7.995 ;
        RECT 866.155 -8.325 866.485 -7.995 ;
        RECT 864.795 -8.325 865.125 -7.995 ;
        RECT 863.435 -8.325 863.765 -7.995 ;
        RECT 862.075 -8.325 862.405 -7.995 ;
        RECT 860.715 -8.325 861.045 -7.995 ;
        RECT 859.355 -8.325 859.685 -7.995 ;
        RECT 857.995 -8.325 858.325 -7.995 ;
        RECT 856.635 -8.325 856.965 -7.995 ;
        RECT 855.275 -8.325 855.605 -7.995 ;
        RECT 853.915 -8.325 854.245 -7.995 ;
        RECT 852.555 -8.325 852.885 -7.995 ;
        RECT 851.195 -8.325 851.525 -7.995 ;
        RECT 849.835 -8.325 850.165 -7.995 ;
        RECT 848.475 -8.325 848.805 -7.995 ;
        RECT 847.115 -8.325 847.445 -7.995 ;
        RECT 845.755 -8.325 846.085 -7.995 ;
        RECT 844.395 -8.325 844.725 -7.995 ;
        RECT 843.035 -8.325 843.365 -7.995 ;
        RECT 841.675 -8.325 842.005 -7.995 ;
        RECT 840.315 -8.325 840.645 -7.995 ;
        RECT 838.955 -8.325 839.285 -7.995 ;
        RECT 837.595 -8.325 837.925 -7.995 ;
        RECT 836.235 -8.325 836.565 -7.995 ;
        RECT 834.875 -8.325 835.205 -7.995 ;
        RECT 833.515 -8.325 833.845 -7.995 ;
        RECT 832.155 -8.325 832.485 -7.995 ;
        RECT 830.795 -8.325 831.125 -7.995 ;
        RECT 829.435 -8.325 829.765 -7.995 ;
        RECT 828.075 -8.325 828.405 -7.995 ;
        RECT 826.715 -8.325 827.045 -7.995 ;
        RECT 825.355 -8.325 825.685 -7.995 ;
        RECT 823.995 -8.325 824.325 -7.995 ;
        RECT 822.635 -8.325 822.965 -7.995 ;
        RECT 821.275 -8.325 821.605 -7.995 ;
        RECT 819.915 -8.325 820.245 -7.995 ;
        RECT 818.555 -8.325 818.885 -7.995 ;
        RECT 817.195 -8.325 817.525 -7.995 ;
        RECT 815.835 -8.325 816.165 -7.995 ;
        RECT 814.475 -8.325 814.805 -7.995 ;
        RECT 813.115 -8.325 813.445 -7.995 ;
        RECT 811.755 -8.325 812.085 -7.995 ;
        RECT 810.395 -8.325 810.725 -7.995 ;
        RECT 809.035 -8.325 809.365 -7.995 ;
        RECT 807.675 -8.325 808.005 -7.995 ;
        RECT 806.315 -8.325 806.645 -7.995 ;
        RECT 804.955 -8.325 805.285 -7.995 ;
        RECT 803.595 -8.325 803.925 -7.995 ;
        RECT 802.235 -8.325 802.565 -7.995 ;
        RECT 800.875 -8.325 801.205 -7.995 ;
        RECT 799.515 -8.325 799.845 -7.995 ;
        RECT 798.155 -8.325 798.485 -7.995 ;
        RECT 796.795 -8.325 797.125 -7.995 ;
        RECT 795.435 -8.325 795.765 -7.995 ;
        RECT 794.075 -8.325 794.405 -7.995 ;
        RECT 792.715 -8.325 793.045 -7.995 ;
        RECT 791.355 -8.325 791.685 -7.995 ;
        RECT 789.995 -8.325 790.325 -7.995 ;
        RECT 788.635 -8.325 788.965 -7.995 ;
        RECT 787.275 -8.325 787.605 -7.995 ;
        RECT 785.915 -8.325 786.245 -7.995 ;
        RECT 784.555 -8.325 784.885 -7.995 ;
        RECT 783.195 -8.325 783.525 -7.995 ;
        RECT 781.835 -8.325 782.165 -7.995 ;
        RECT 780.475 -8.325 780.805 -7.995 ;
        RECT 779.115 -8.325 779.445 -7.995 ;
        RECT 777.755 -8.325 778.085 -7.995 ;
        RECT 776.395 -8.325 776.725 -7.995 ;
        RECT 775.035 -8.325 775.365 -7.995 ;
        RECT 773.675 -8.325 774.005 -7.995 ;
        RECT 772.315 -8.325 772.645 -7.995 ;
        RECT 770.955 -8.325 771.285 -7.995 ;
        RECT 769.595 -8.325 769.925 -7.995 ;
        RECT 768.235 -8.325 768.565 -7.995 ;
        RECT 766.875 -8.325 767.205 -7.995 ;
        RECT 765.515 -8.325 765.845 -7.995 ;
        RECT 764.155 -8.325 764.485 -7.995 ;
        RECT 762.795 -8.325 763.125 -7.995 ;
        RECT 761.435 -8.325 761.765 -7.995 ;
        RECT 760.075 -8.325 760.405 -7.995 ;
        RECT 758.715 -8.325 759.045 -7.995 ;
        RECT 757.355 -8.325 757.685 -7.995 ;
        RECT 755.995 -8.325 756.325 -7.995 ;
        RECT 754.635 -8.325 754.965 -7.995 ;
        RECT 753.275 -8.325 753.605 -7.995 ;
        RECT 751.915 -8.325 752.245 -7.995 ;
        RECT 750.555 -8.325 750.885 -7.995 ;
        RECT 749.195 -8.325 749.525 -7.995 ;
        RECT 747.835 -8.325 748.165 -7.995 ;
        RECT 746.475 -8.325 746.805 -7.995 ;
        RECT 745.115 -8.325 745.445 -7.995 ;
        RECT 743.755 -8.325 744.085 -7.995 ;
        RECT 742.395 -8.325 742.725 -7.995 ;
        RECT 741.035 -8.325 741.365 -7.995 ;
        RECT 739.675 -8.325 740.005 -7.995 ;
        RECT 738.315 -8.325 738.645 -7.995 ;
        RECT 736.955 -8.325 737.285 -7.995 ;
        RECT 735.595 -8.325 735.925 -7.995 ;
        RECT 734.235 -8.325 734.565 -7.995 ;
        RECT 732.875 -8.325 733.205 -7.995 ;
        RECT 731.515 -8.325 731.845 -7.995 ;
        RECT 730.155 -8.325 730.485 -7.995 ;
        RECT 728.795 -8.325 729.125 -7.995 ;
        RECT 727.435 -8.325 727.765 -7.995 ;
        RECT 726.075 -8.325 726.405 -7.995 ;
        RECT 724.715 -8.325 725.045 -7.995 ;
        RECT 723.355 -8.325 723.685 -7.995 ;
        RECT 721.995 -8.325 722.325 -7.995 ;
        RECT 720.635 -8.325 720.965 -7.995 ;
        RECT 719.275 -8.325 719.605 -7.995 ;
        RECT 717.915 -8.325 718.245 -7.995 ;
        RECT 716.555 -8.325 716.885 -7.995 ;
        RECT 715.195 -8.325 715.525 -7.995 ;
        RECT 713.835 -8.325 714.165 -7.995 ;
        RECT 712.475 -8.325 712.805 -7.995 ;
        RECT 711.115 -8.325 711.445 -7.995 ;
        RECT 709.755 -8.325 710.085 -7.995 ;
        RECT 708.395 -8.325 708.725 -7.995 ;
        RECT 707.035 -8.325 707.365 -7.995 ;
        RECT 705.675 -8.325 706.005 -7.995 ;
        RECT 704.315 -8.325 704.645 -7.995 ;
        RECT 702.955 -8.325 703.285 -7.995 ;
        RECT 701.595 -8.325 701.925 -7.995 ;
        RECT 700.235 -8.325 700.565 -7.995 ;
        RECT 698.875 -8.325 699.205 -7.995 ;
        RECT 697.515 -8.325 697.845 -7.995 ;
        RECT 696.155 -8.325 696.485 -7.995 ;
        RECT 694.795 -8.325 695.125 -7.995 ;
        RECT 693.435 -8.325 693.765 -7.995 ;
        RECT 692.075 -8.325 692.405 -7.995 ;
        RECT 690.715 -8.325 691.045 -7.995 ;
        RECT 689.355 -8.325 689.685 -7.995 ;
        RECT 687.995 -8.325 688.325 -7.995 ;
        RECT 686.635 -8.325 686.965 -7.995 ;
        RECT 685.275 -8.325 685.605 -7.995 ;
        RECT 683.915 -8.325 684.245 -7.995 ;
        RECT 682.555 -8.325 682.885 -7.995 ;
        RECT 681.195 -8.325 681.525 -7.995 ;
        RECT 679.835 -8.325 680.165 -7.995 ;
        RECT 678.475 -8.325 678.805 -7.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -4.24 678.475 -3.92 ;
        RECT 677.115 -4.245 677.445 -3.915 ;
        RECT 675.755 -4.245 676.085 -3.915 ;
        RECT 674.395 -4.245 674.725 -3.915 ;
        RECT 673.035 -4.245 673.365 -3.915 ;
        RECT 671.675 -4.245 672.005 -3.915 ;
        RECT 670.315 -4.245 670.645 -3.915 ;
        RECT 668.955 -4.245 669.285 -3.915 ;
        RECT 667.595 -4.245 667.925 -3.915 ;
        RECT 666.235 -4.245 666.565 -3.915 ;
        RECT 664.875 -4.245 665.205 -3.915 ;
        RECT 663.515 -4.245 663.845 -3.915 ;
        RECT 662.155 -4.245 662.485 -3.915 ;
        RECT 660.795 -4.245 661.125 -3.915 ;
        RECT 659.435 -4.245 659.765 -3.915 ;
        RECT 658.075 -4.245 658.405 -3.915 ;
        RECT 656.715 -4.245 657.045 -3.915 ;
        RECT 655.355 -4.245 655.685 -3.915 ;
        RECT 653.995 -4.245 654.325 -3.915 ;
        RECT 652.635 -4.245 652.965 -3.915 ;
        RECT 651.275 -4.245 651.605 -3.915 ;
        RECT 649.915 -4.245 650.245 -3.915 ;
        RECT 648.555 -4.245 648.885 -3.915 ;
        RECT 647.195 -4.245 647.525 -3.915 ;
        RECT 645.835 -4.245 646.165 -3.915 ;
        RECT 644.475 -4.245 644.805 -3.915 ;
        RECT 643.115 -4.245 643.445 -3.915 ;
        RECT 641.755 -4.245 642.085 -3.915 ;
        RECT 640.395 -4.245 640.725 -3.915 ;
        RECT 639.035 -4.245 639.365 -3.915 ;
        RECT 637.675 -4.245 638.005 -3.915 ;
        RECT 636.315 -4.245 636.645 -3.915 ;
        RECT 634.955 -4.245 635.285 -3.915 ;
        RECT 633.595 -4.245 633.925 -3.915 ;
        RECT 632.235 -4.245 632.565 -3.915 ;
        RECT 630.875 -4.245 631.205 -3.915 ;
        RECT 629.515 -4.245 629.845 -3.915 ;
        RECT 628.155 -4.245 628.485 -3.915 ;
        RECT 626.795 -4.245 627.125 -3.915 ;
        RECT 625.435 -4.245 625.765 -3.915 ;
        RECT 624.075 -4.245 624.405 -3.915 ;
        RECT 622.715 -4.245 623.045 -3.915 ;
        RECT 621.355 -4.245 621.685 -3.915 ;
        RECT 619.995 -4.245 620.325 -3.915 ;
        RECT 618.635 -4.245 618.965 -3.915 ;
        RECT 617.275 -4.245 617.605 -3.915 ;
        RECT 615.915 -4.245 616.245 -3.915 ;
        RECT 614.555 -4.245 614.885 -3.915 ;
        RECT 613.195 -4.245 613.525 -3.915 ;
        RECT 611.835 -4.245 612.165 -3.915 ;
        RECT 610.475 -4.245 610.805 -3.915 ;
        RECT 609.115 -4.245 609.445 -3.915 ;
        RECT 607.755 -4.245 608.085 -3.915 ;
        RECT 606.395 -4.245 606.725 -3.915 ;
        RECT 605.035 -4.245 605.365 -3.915 ;
        RECT 603.675 -4.245 604.005 -3.915 ;
        RECT 602.315 -4.245 602.645 -3.915 ;
        RECT 600.955 -4.245 601.285 -3.915 ;
        RECT 599.595 -4.245 599.925 -3.915 ;
        RECT 598.235 -4.245 598.565 -3.915 ;
        RECT 596.875 -4.245 597.205 -3.915 ;
        RECT 595.515 -4.245 595.845 -3.915 ;
        RECT 594.155 -4.245 594.485 -3.915 ;
        RECT 592.795 -4.245 593.125 -3.915 ;
        RECT 591.435 -4.245 591.765 -3.915 ;
        RECT 590.075 -4.245 590.405 -3.915 ;
        RECT 588.715 -4.245 589.045 -3.915 ;
        RECT 587.355 -4.245 587.685 -3.915 ;
        RECT 585.995 -4.245 586.325 -3.915 ;
        RECT 584.635 -4.245 584.965 -3.915 ;
        RECT 583.275 -4.245 583.605 -3.915 ;
        RECT 581.915 -4.245 582.245 -3.915 ;
        RECT 580.555 -4.245 580.885 -3.915 ;
        RECT 579.195 -4.245 579.525 -3.915 ;
        RECT 577.835 -4.245 578.165 -3.915 ;
        RECT 576.475 -4.245 576.805 -3.915 ;
        RECT 575.115 -4.245 575.445 -3.915 ;
        RECT 573.755 -4.245 574.085 -3.915 ;
        RECT 572.395 -4.245 572.725 -3.915 ;
        RECT 571.035 -4.245 571.365 -3.915 ;
        RECT 569.675 -4.245 570.005 -3.915 ;
        RECT 568.315 -4.245 568.645 -3.915 ;
        RECT 566.955 -4.245 567.285 -3.915 ;
        RECT 565.595 -4.245 565.925 -3.915 ;
        RECT 564.235 -4.245 564.565 -3.915 ;
        RECT 562.875 -4.245 563.205 -3.915 ;
        RECT 561.515 -4.245 561.845 -3.915 ;
        RECT 560.155 -4.245 560.485 -3.915 ;
        RECT 558.795 -4.245 559.125 -3.915 ;
        RECT 557.435 -4.245 557.765 -3.915 ;
        RECT 556.075 -4.245 556.405 -3.915 ;
        RECT 554.715 -4.245 555.045 -3.915 ;
        RECT 553.355 -4.245 553.685 -3.915 ;
        RECT 551.995 -4.245 552.325 -3.915 ;
        RECT 550.635 -4.245 550.965 -3.915 ;
        RECT 549.275 -4.245 549.605 -3.915 ;
        RECT 547.915 -4.245 548.245 -3.915 ;
        RECT 546.555 -4.245 546.885 -3.915 ;
        RECT 545.195 -4.245 545.525 -3.915 ;
        RECT 543.835 -4.245 544.165 -3.915 ;
        RECT 542.475 -4.245 542.805 -3.915 ;
        RECT 541.115 -4.245 541.445 -3.915 ;
        RECT 539.755 -4.245 540.085 -3.915 ;
        RECT 538.395 -4.245 538.725 -3.915 ;
        RECT 537.035 -4.245 537.365 -3.915 ;
        RECT 535.675 -4.245 536.005 -3.915 ;
        RECT 534.315 -4.245 534.645 -3.915 ;
        RECT 532.955 -4.245 533.285 -3.915 ;
        RECT 531.595 -4.245 531.925 -3.915 ;
        RECT 530.235 -4.245 530.565 -3.915 ;
        RECT 528.875 -4.245 529.205 -3.915 ;
        RECT 527.515 -4.245 527.845 -3.915 ;
        RECT 526.155 -4.245 526.485 -3.915 ;
        RECT 524.795 -4.245 525.125 -3.915 ;
        RECT 523.435 -4.245 523.765 -3.915 ;
        RECT 522.075 -4.245 522.405 -3.915 ;
        RECT 520.715 -4.245 521.045 -3.915 ;
        RECT 519.355 -4.245 519.685 -3.915 ;
        RECT 517.995 -4.245 518.325 -3.915 ;
        RECT 516.635 -4.245 516.965 -3.915 ;
        RECT 515.275 -4.245 515.605 -3.915 ;
        RECT 513.915 -4.245 514.245 -3.915 ;
        RECT 512.555 -4.245 512.885 -3.915 ;
        RECT 511.195 -4.245 511.525 -3.915 ;
        RECT 509.835 -4.245 510.165 -3.915 ;
        RECT 508.475 -4.245 508.805 -3.915 ;
        RECT 507.115 -4.245 507.445 -3.915 ;
        RECT 505.755 -4.245 506.085 -3.915 ;
        RECT 504.395 -4.245 504.725 -3.915 ;
        RECT 503.035 -4.245 503.365 -3.915 ;
        RECT 501.675 -4.245 502.005 -3.915 ;
        RECT 500.315 -4.245 500.645 -3.915 ;
        RECT 498.955 -4.245 499.285 -3.915 ;
        RECT 497.595 -4.245 497.925 -3.915 ;
        RECT 496.235 -4.245 496.565 -3.915 ;
        RECT 494.875 -4.245 495.205 -3.915 ;
        RECT 493.515 -4.245 493.845 -3.915 ;
        RECT 492.155 -4.245 492.485 -3.915 ;
        RECT 490.795 -4.245 491.125 -3.915 ;
        RECT 489.435 -4.245 489.765 -3.915 ;
        RECT 488.075 -4.245 488.405 -3.915 ;
        RECT 486.715 -4.245 487.045 -3.915 ;
        RECT 485.355 -4.245 485.685 -3.915 ;
        RECT 483.995 -4.245 484.325 -3.915 ;
        RECT 482.635 -4.245 482.965 -3.915 ;
        RECT 481.275 -4.245 481.605 -3.915 ;
        RECT 479.915 -4.245 480.245 -3.915 ;
        RECT 478.555 -4.245 478.885 -3.915 ;
        RECT 477.195 -4.245 477.525 -3.915 ;
        RECT 475.835 -4.245 476.165 -3.915 ;
        RECT 474.475 -4.245 474.805 -3.915 ;
        RECT 473.115 -4.245 473.445 -3.915 ;
        RECT 471.755 -4.245 472.085 -3.915 ;
        RECT 470.395 -4.245 470.725 -3.915 ;
        RECT 469.035 -4.245 469.365 -3.915 ;
        RECT 467.675 -4.245 468.005 -3.915 ;
        RECT 466.315 -4.245 466.645 -3.915 ;
        RECT 464.955 -4.245 465.285 -3.915 ;
        RECT 463.595 -4.245 463.925 -3.915 ;
        RECT 462.235 -4.245 462.565 -3.915 ;
        RECT 460.875 -4.245 461.205 -3.915 ;
        RECT 459.515 -4.245 459.845 -3.915 ;
        RECT 458.155 -4.245 458.485 -3.915 ;
        RECT 456.795 -4.245 457.125 -3.915 ;
        RECT 455.435 -4.245 455.765 -3.915 ;
        RECT 454.075 -4.245 454.405 -3.915 ;
        RECT 452.715 -4.245 453.045 -3.915 ;
        RECT 451.355 -4.245 451.685 -3.915 ;
        RECT 449.995 -4.245 450.325 -3.915 ;
        RECT 448.635 -4.245 448.965 -3.915 ;
        RECT 447.275 -4.245 447.605 -3.915 ;
        RECT 445.915 -4.245 446.245 -3.915 ;
        RECT 444.555 -4.245 444.885 -3.915 ;
        RECT 443.195 -4.245 443.525 -3.915 ;
        RECT 441.835 -4.245 442.165 -3.915 ;
        RECT 440.475 -4.245 440.805 -3.915 ;
        RECT 439.115 -4.245 439.445 -3.915 ;
        RECT 437.755 -4.245 438.085 -3.915 ;
        RECT 436.395 -4.245 436.725 -3.915 ;
        RECT 435.035 -4.245 435.365 -3.915 ;
        RECT 433.675 -4.245 434.005 -3.915 ;
        RECT 432.315 -4.245 432.645 -3.915 ;
        RECT 430.955 -4.245 431.285 -3.915 ;
        RECT 429.595 -4.245 429.925 -3.915 ;
        RECT 428.235 -4.245 428.565 -3.915 ;
        RECT 426.875 -4.245 427.205 -3.915 ;
        RECT 425.515 -4.245 425.845 -3.915 ;
        RECT 424.155 -4.245 424.485 -3.915 ;
        RECT 422.795 -4.245 423.125 -3.915 ;
        RECT 421.435 -4.245 421.765 -3.915 ;
        RECT 420.075 -4.245 420.405 -3.915 ;
        RECT 418.715 -4.245 419.045 -3.915 ;
        RECT 417.355 -4.245 417.685 -3.915 ;
        RECT 415.995 -4.245 416.325 -3.915 ;
        RECT 414.635 -4.245 414.965 -3.915 ;
        RECT 413.275 -4.245 413.605 -3.915 ;
        RECT 411.915 -4.245 412.245 -3.915 ;
        RECT 410.555 -4.245 410.885 -3.915 ;
        RECT 409.195 -4.245 409.525 -3.915 ;
        RECT 407.835 -4.245 408.165 -3.915 ;
        RECT 406.475 -4.245 406.805 -3.915 ;
        RECT 405.115 -4.245 405.445 -3.915 ;
        RECT 403.755 -4.245 404.085 -3.915 ;
        RECT 402.395 -4.245 402.725 -3.915 ;
        RECT 401.035 -4.245 401.365 -3.915 ;
        RECT 399.675 -4.245 400.005 -3.915 ;
        RECT 398.315 -4.245 398.645 -3.915 ;
        RECT 396.955 -4.245 397.285 -3.915 ;
        RECT 395.595 -4.245 395.925 -3.915 ;
        RECT 394.235 -4.245 394.565 -3.915 ;
        RECT 392.875 -4.245 393.205 -3.915 ;
        RECT 391.515 -4.245 391.845 -3.915 ;
        RECT 390.155 -4.245 390.485 -3.915 ;
        RECT 388.795 -4.245 389.125 -3.915 ;
        RECT 387.435 -4.245 387.765 -3.915 ;
        RECT 386.075 -4.245 386.405 -3.915 ;
        RECT 384.715 -4.245 385.045 -3.915 ;
        RECT 383.355 -4.245 383.685 -3.915 ;
        RECT 381.995 -4.245 382.325 -3.915 ;
        RECT 380.635 -4.245 380.965 -3.915 ;
        RECT 379.275 -4.245 379.605 -3.915 ;
        RECT 377.915 -4.245 378.245 -3.915 ;
        RECT 376.555 -4.245 376.885 -3.915 ;
        RECT 375.195 -4.245 375.525 -3.915 ;
        RECT 373.835 -4.245 374.165 -3.915 ;
        RECT 372.475 -4.245 372.805 -3.915 ;
        RECT 371.115 -4.245 371.445 -3.915 ;
        RECT 369.755 -4.245 370.085 -3.915 ;
        RECT 368.395 -4.245 368.725 -3.915 ;
        RECT 367.035 -4.245 367.365 -3.915 ;
        RECT 365.675 -4.245 366.005 -3.915 ;
        RECT 364.315 -4.245 364.645 -3.915 ;
        RECT 362.955 -4.245 363.285 -3.915 ;
        RECT 361.595 -4.245 361.925 -3.915 ;
        RECT 360.235 -4.245 360.565 -3.915 ;
        RECT 358.875 -4.245 359.205 -3.915 ;
        RECT 357.515 -4.245 357.845 -3.915 ;
        RECT 356.155 -4.245 356.485 -3.915 ;
        RECT 354.795 -4.245 355.125 -3.915 ;
        RECT 353.435 -4.245 353.765 -3.915 ;
        RECT 352.075 -4.245 352.405 -3.915 ;
        RECT 350.715 -4.245 351.045 -3.915 ;
        RECT 349.355 -4.245 349.685 -3.915 ;
        RECT 347.995 -4.245 348.325 -3.915 ;
        RECT 346.635 -4.245 346.965 -3.915 ;
        RECT 345.275 -4.245 345.605 -3.915 ;
        RECT 343.915 -4.245 344.245 -3.915 ;
        RECT 342.555 -4.245 342.885 -3.915 ;
        RECT 341.195 -4.245 341.525 -3.915 ;
        RECT 339.835 -4.245 340.165 -3.915 ;
        RECT 338.475 -4.245 338.805 -3.915 ;
        RECT 337.115 -4.245 337.445 -3.915 ;
        RECT 335.755 -4.245 336.085 -3.915 ;
        RECT 334.395 -4.245 334.725 -3.915 ;
        RECT 333.035 -4.245 333.365 -3.915 ;
        RECT 331.675 -4.245 332.005 -3.915 ;
        RECT 330.315 -4.245 330.645 -3.915 ;
        RECT 328.955 -4.245 329.285 -3.915 ;
        RECT 327.595 -4.245 327.925 -3.915 ;
        RECT 326.235 -4.245 326.565 -3.915 ;
        RECT 324.875 -4.245 325.205 -3.915 ;
        RECT 323.515 -4.245 323.845 -3.915 ;
        RECT 322.155 -4.245 322.485 -3.915 ;
        RECT 320.795 -4.245 321.125 -3.915 ;
        RECT 319.435 -4.245 319.765 -3.915 ;
        RECT 318.075 -4.245 318.405 -3.915 ;
        RECT 316.715 -4.245 317.045 -3.915 ;
        RECT 315.355 -4.245 315.685 -3.915 ;
        RECT 313.995 -4.245 314.325 -3.915 ;
        RECT 312.635 -4.245 312.965 -3.915 ;
        RECT 311.275 -4.245 311.605 -3.915 ;
        RECT 309.915 -4.245 310.245 -3.915 ;
        RECT 308.555 -4.245 308.885 -3.915 ;
        RECT 307.195 -4.245 307.525 -3.915 ;
        RECT 305.835 -4.245 306.165 -3.915 ;
        RECT 304.475 -4.245 304.805 -3.915 ;
        RECT 303.115 -4.245 303.445 -3.915 ;
        RECT 301.755 -4.245 302.085 -3.915 ;
        RECT 300.395 -4.245 300.725 -3.915 ;
        RECT 299.035 -4.245 299.365 -3.915 ;
        RECT 297.675 -4.245 298.005 -3.915 ;
        RECT 296.315 -4.245 296.645 -3.915 ;
        RECT 294.955 -4.245 295.285 -3.915 ;
        RECT 293.595 -4.245 293.925 -3.915 ;
        RECT 292.235 -4.245 292.565 -3.915 ;
        RECT 290.875 -4.245 291.205 -3.915 ;
        RECT 289.515 -4.245 289.845 -3.915 ;
        RECT 288.155 -4.245 288.485 -3.915 ;
        RECT 286.795 -4.245 287.125 -3.915 ;
        RECT 285.435 -4.245 285.765 -3.915 ;
        RECT 284.075 -4.245 284.405 -3.915 ;
        RECT 282.715 -4.245 283.045 -3.915 ;
        RECT 281.355 -4.245 281.685 -3.915 ;
        RECT 279.995 -4.245 280.325 -3.915 ;
        RECT 278.635 -4.245 278.965 -3.915 ;
        RECT 277.275 -4.245 277.605 -3.915 ;
        RECT 275.915 -4.245 276.245 -3.915 ;
        RECT 274.555 -4.245 274.885 -3.915 ;
        RECT 273.195 -4.245 273.525 -3.915 ;
        RECT 271.835 -4.245 272.165 -3.915 ;
        RECT 270.475 -4.245 270.805 -3.915 ;
        RECT 269.115 -4.245 269.445 -3.915 ;
        RECT 267.755 -4.245 268.085 -3.915 ;
        RECT 266.395 -4.245 266.725 -3.915 ;
        RECT 265.035 -4.245 265.365 -3.915 ;
        RECT 263.675 -4.245 264.005 -3.915 ;
        RECT 262.315 -4.245 262.645 -3.915 ;
        RECT 260.955 -4.245 261.285 -3.915 ;
        RECT 259.595 -4.245 259.925 -3.915 ;
        RECT 258.235 -4.245 258.565 -3.915 ;
        RECT 256.875 -4.245 257.205 -3.915 ;
        RECT 255.515 -4.245 255.845 -3.915 ;
        RECT 254.155 -4.245 254.485 -3.915 ;
        RECT 252.795 -4.245 253.125 -3.915 ;
        RECT 251.435 -4.245 251.765 -3.915 ;
        RECT 250.075 -4.245 250.405 -3.915 ;
        RECT 248.715 -4.245 249.045 -3.915 ;
        RECT 247.355 -4.245 247.685 -3.915 ;
        RECT 245.995 -4.245 246.325 -3.915 ;
        RECT 244.635 -4.245 244.965 -3.915 ;
        RECT 243.275 -4.245 243.605 -3.915 ;
        RECT 241.915 -4.245 242.245 -3.915 ;
        RECT 240.555 -4.245 240.885 -3.915 ;
        RECT 239.195 -4.245 239.525 -3.915 ;
        RECT 237.835 -4.245 238.165 -3.915 ;
        RECT 236.475 -4.245 236.805 -3.915 ;
        RECT 235.115 -4.245 235.445 -3.915 ;
        RECT 233.755 -4.245 234.085 -3.915 ;
        RECT 232.395 -4.245 232.725 -3.915 ;
        RECT 231.035 -4.245 231.365 -3.915 ;
        RECT 229.675 -4.245 230.005 -3.915 ;
        RECT 228.315 -4.245 228.645 -3.915 ;
        RECT 226.955 -4.245 227.285 -3.915 ;
        RECT 225.595 -4.245 225.925 -3.915 ;
        RECT 224.235 -4.245 224.565 -3.915 ;
        RECT 222.875 -4.245 223.205 -3.915 ;
        RECT 221.515 -4.245 221.845 -3.915 ;
        RECT 220.155 -4.245 220.485 -3.915 ;
        RECT 218.795 -4.245 219.125 -3.915 ;
        RECT 217.435 -4.245 217.765 -3.915 ;
        RECT 216.075 -4.245 216.405 -3.915 ;
        RECT 214.715 -4.245 215.045 -3.915 ;
        RECT 213.355 -4.245 213.685 -3.915 ;
        RECT 211.995 -4.245 212.325 -3.915 ;
        RECT 210.635 -4.245 210.965 -3.915 ;
        RECT 209.275 -4.245 209.605 -3.915 ;
        RECT 207.915 -4.245 208.245 -3.915 ;
        RECT 206.555 -4.245 206.885 -3.915 ;
        RECT 205.195 -4.245 205.525 -3.915 ;
        RECT 203.835 -4.245 204.165 -3.915 ;
        RECT 202.475 -4.245 202.805 -3.915 ;
        RECT 201.115 -4.245 201.445 -3.915 ;
        RECT 199.755 -4.245 200.085 -3.915 ;
        RECT 198.395 -4.245 198.725 -3.915 ;
        RECT 197.035 -4.245 197.365 -3.915 ;
        RECT 195.675 -4.245 196.005 -3.915 ;
        RECT 194.315 -4.245 194.645 -3.915 ;
        RECT 192.955 -4.245 193.285 -3.915 ;
        RECT 191.595 -4.245 191.925 -3.915 ;
        RECT 190.235 -4.245 190.565 -3.915 ;
        RECT 188.875 -4.245 189.205 -3.915 ;
        RECT 187.515 -4.245 187.845 -3.915 ;
        RECT 186.155 -4.245 186.485 -3.915 ;
        RECT 184.795 -4.245 185.125 -3.915 ;
        RECT 183.435 -4.245 183.765 -3.915 ;
        RECT 182.075 -4.245 182.405 -3.915 ;
        RECT 180.715 -4.245 181.045 -3.915 ;
        RECT 179.355 -4.245 179.685 -3.915 ;
        RECT 177.995 -4.245 178.325 -3.915 ;
        RECT 176.635 -4.245 176.965 -3.915 ;
        RECT 175.275 -4.245 175.605 -3.915 ;
        RECT 173.915 -4.245 174.245 -3.915 ;
        RECT 172.555 -4.245 172.885 -3.915 ;
        RECT 171.195 -4.245 171.525 -3.915 ;
        RECT 169.835 -4.245 170.165 -3.915 ;
        RECT 168.475 -4.245 168.805 -3.915 ;
        RECT 167.115 -4.245 167.445 -3.915 ;
        RECT 165.755 -4.245 166.085 -3.915 ;
        RECT 164.395 -4.245 164.725 -3.915 ;
        RECT 163.035 -4.245 163.365 -3.915 ;
        RECT 161.675 -4.245 162.005 -3.915 ;
        RECT 160.315 -4.245 160.645 -3.915 ;
        RECT 158.955 -4.245 159.285 -3.915 ;
        RECT 157.595 -4.245 157.925 -3.915 ;
        RECT 156.235 -4.245 156.565 -3.915 ;
        RECT 154.875 -4.245 155.205 -3.915 ;
        RECT 153.515 -4.245 153.845 -3.915 ;
        RECT 152.155 -4.245 152.485 -3.915 ;
        RECT 150.795 -4.245 151.125 -3.915 ;
        RECT 149.435 -4.245 149.765 -3.915 ;
        RECT 148.075 -4.245 148.405 -3.915 ;
        RECT 146.715 -4.245 147.045 -3.915 ;
        RECT 145.355 -4.245 145.685 -3.915 ;
        RECT 143.995 -4.245 144.325 -3.915 ;
        RECT 142.635 -4.245 142.965 -3.915 ;
        RECT 141.275 -4.245 141.605 -3.915 ;
        RECT 139.915 -4.245 140.245 -3.915 ;
        RECT 138.555 -4.245 138.885 -3.915 ;
        RECT 137.195 -4.245 137.525 -3.915 ;
        RECT 135.835 -4.245 136.165 -3.915 ;
        RECT 134.475 -4.245 134.805 -3.915 ;
        RECT 133.115 -4.245 133.445 -3.915 ;
        RECT 131.755 -4.245 132.085 -3.915 ;
        RECT 130.395 -4.245 130.725 -3.915 ;
        RECT 129.035 -4.245 129.365 -3.915 ;
        RECT 127.675 -4.245 128.005 -3.915 ;
        RECT 126.315 -4.245 126.645 -3.915 ;
        RECT 124.955 -4.245 125.285 -3.915 ;
        RECT 123.595 -4.245 123.925 -3.915 ;
        RECT 122.235 -4.245 122.565 -3.915 ;
        RECT 120.875 -4.245 121.205 -3.915 ;
        RECT 119.515 -4.245 119.845 -3.915 ;
        RECT 118.155 -4.245 118.485 -3.915 ;
        RECT 116.795 -4.245 117.125 -3.915 ;
        RECT 115.435 -4.245 115.765 -3.915 ;
        RECT 114.075 -4.245 114.405 -3.915 ;
        RECT 112.715 -4.245 113.045 -3.915 ;
        RECT 111.355 -4.245 111.685 -3.915 ;
        RECT 109.995 -4.245 110.325 -3.915 ;
        RECT 108.635 -4.245 108.965 -3.915 ;
        RECT 107.275 -4.245 107.605 -3.915 ;
        RECT 105.915 -4.245 106.245 -3.915 ;
        RECT 104.555 -4.245 104.885 -3.915 ;
        RECT 103.195 -4.245 103.525 -3.915 ;
        RECT 101.835 -4.245 102.165 -3.915 ;
        RECT 100.475 -4.245 100.805 -3.915 ;
        RECT 99.115 -4.245 99.445 -3.915 ;
        RECT 97.755 -4.245 98.085 -3.915 ;
        RECT 96.395 -4.245 96.725 -3.915 ;
        RECT 95.035 -4.245 95.365 -3.915 ;
        RECT 93.675 -4.245 94.005 -3.915 ;
        RECT 92.315 -4.245 92.645 -3.915 ;
        RECT 90.955 -4.245 91.285 -3.915 ;
        RECT 89.595 -4.245 89.925 -3.915 ;
        RECT 88.235 -4.245 88.565 -3.915 ;
        RECT 86.875 -4.245 87.205 -3.915 ;
        RECT 85.515 -4.245 85.845 -3.915 ;
        RECT 84.155 -4.245 84.485 -3.915 ;
        RECT 82.795 -4.245 83.125 -3.915 ;
        RECT 81.435 -4.245 81.765 -3.915 ;
        RECT 80.075 -4.245 80.405 -3.915 ;
        RECT 78.715 -4.245 79.045 -3.915 ;
        RECT 77.355 -4.245 77.685 -3.915 ;
        RECT 75.995 -4.245 76.325 -3.915 ;
        RECT 74.635 -4.245 74.965 -3.915 ;
        RECT 73.275 -4.245 73.605 -3.915 ;
        RECT 71.915 -4.245 72.245 -3.915 ;
        RECT 70.555 -4.245 70.885 -3.915 ;
        RECT 69.195 -4.245 69.525 -3.915 ;
        RECT 67.835 -4.245 68.165 -3.915 ;
        RECT 66.475 -4.245 66.805 -3.915 ;
        RECT 65.115 -4.245 65.445 -3.915 ;
        RECT 63.755 -4.245 64.085 -3.915 ;
        RECT 62.395 -4.245 62.725 -3.915 ;
        RECT 61.035 -4.245 61.365 -3.915 ;
        RECT 59.675 -4.245 60.005 -3.915 ;
        RECT 58.315 -4.245 58.645 -3.915 ;
        RECT 56.955 -4.245 57.285 -3.915 ;
        RECT 55.595 -4.245 55.925 -3.915 ;
        RECT 54.235 -4.245 54.565 -3.915 ;
        RECT 52.875 -4.245 53.205 -3.915 ;
        RECT 51.515 -4.245 51.845 -3.915 ;
        RECT 50.155 -4.245 50.485 -3.915 ;
        RECT 48.795 -4.245 49.125 -3.915 ;
        RECT 47.435 -4.245 47.765 -3.915 ;
        RECT 46.075 -4.245 46.405 -3.915 ;
        RECT 44.715 -4.245 45.045 -3.915 ;
        RECT 43.355 -4.245 43.685 -3.915 ;
        RECT 41.995 -4.245 42.325 -3.915 ;
        RECT 40.635 -4.245 40.965 -3.915 ;
        RECT 39.275 -4.245 39.605 -3.915 ;
        RECT 37.915 -4.245 38.245 -3.915 ;
        RECT 36.555 -4.245 36.885 -3.915 ;
        RECT 35.195 -4.245 35.525 -3.915 ;
        RECT 33.835 -4.245 34.165 -3.915 ;
        RECT 32.475 -4.245 32.805 -3.915 ;
        RECT 31.115 -4.245 31.445 -3.915 ;
        RECT 29.755 -4.245 30.085 -3.915 ;
        RECT 28.395 -4.245 28.725 -3.915 ;
        RECT 27.035 -4.245 27.365 -3.915 ;
        RECT 25.675 -4.245 26.005 -3.915 ;
        RECT 24.315 -4.245 24.645 -3.915 ;
        RECT 22.955 -4.245 23.285 -3.915 ;
        RECT 21.595 -4.245 21.925 -3.915 ;
        RECT 20.235 -4.245 20.565 -3.915 ;
        RECT 18.875 -4.245 19.205 -3.915 ;
        RECT 17.515 -4.245 17.845 -3.915 ;
        RECT 16.155 -4.245 16.485 -3.915 ;
        RECT 14.795 -4.245 15.125 -3.915 ;
        RECT 13.435 -4.245 13.765 -3.915 ;
        RECT 12.075 -4.245 12.405 -3.915 ;
        RECT 10.715 -4.245 11.045 -3.915 ;
        RECT 9.355 -4.245 9.685 -3.915 ;
        RECT 7.995 -4.245 8.325 -3.915 ;
        RECT 6.635 -4.245 6.965 -3.915 ;
        RECT 5.275 -4.245 5.605 -3.915 ;
        RECT 3.915 -4.245 4.245 -3.915 ;
        RECT 2.555 -4.245 2.885 -3.915 ;
        RECT 1.195 -4.245 1.525 -3.915 ;
        RECT -0.165 -4.245 0.165 -3.915 ;
        RECT -1.525 -4.245 -1.195 -3.915 ;
        RECT 874.315 -4.245 874.645 -3.915 ;
        RECT 872.955 -4.245 873.285 -3.915 ;
        RECT 871.595 -4.245 871.925 -3.915 ;
        RECT 870.235 -4.245 870.565 -3.915 ;
        RECT 868.875 -4.245 869.205 -3.915 ;
        RECT 867.515 -4.245 867.845 -3.915 ;
        RECT 866.155 -4.245 866.485 -3.915 ;
        RECT 864.795 -4.245 865.125 -3.915 ;
        RECT 863.435 -4.245 863.765 -3.915 ;
        RECT 862.075 -4.245 862.405 -3.915 ;
        RECT 860.715 -4.245 861.045 -3.915 ;
        RECT 859.355 -4.245 859.685 -3.915 ;
        RECT 857.995 -4.245 858.325 -3.915 ;
        RECT 856.635 -4.245 856.965 -3.915 ;
        RECT 855.275 -4.245 855.605 -3.915 ;
        RECT 853.915 -4.245 854.245 -3.915 ;
        RECT 852.555 -4.245 852.885 -3.915 ;
        RECT 851.195 -4.245 851.525 -3.915 ;
        RECT 849.835 -4.245 850.165 -3.915 ;
        RECT 848.475 -4.245 848.805 -3.915 ;
        RECT 847.115 -4.245 847.445 -3.915 ;
        RECT 845.755 -4.245 846.085 -3.915 ;
        RECT 844.395 -4.245 844.725 -3.915 ;
        RECT 843.035 -4.245 843.365 -3.915 ;
        RECT 841.675 -4.245 842.005 -3.915 ;
        RECT 840.315 -4.245 840.645 -3.915 ;
        RECT 838.955 -4.245 839.285 -3.915 ;
        RECT 837.595 -4.245 837.925 -3.915 ;
        RECT 836.235 -4.245 836.565 -3.915 ;
        RECT 834.875 -4.245 835.205 -3.915 ;
        RECT 833.515 -4.245 833.845 -3.915 ;
        RECT 832.155 -4.245 832.485 -3.915 ;
        RECT 830.795 -4.245 831.125 -3.915 ;
        RECT 829.435 -4.245 829.765 -3.915 ;
        RECT 828.075 -4.245 828.405 -3.915 ;
        RECT 826.715 -4.245 827.045 -3.915 ;
        RECT 825.355 -4.245 825.685 -3.915 ;
        RECT 823.995 -4.245 824.325 -3.915 ;
        RECT 822.635 -4.245 822.965 -3.915 ;
        RECT 821.275 -4.245 821.605 -3.915 ;
        RECT 819.915 -4.245 820.245 -3.915 ;
        RECT 818.555 -4.245 818.885 -3.915 ;
        RECT 817.195 -4.245 817.525 -3.915 ;
        RECT 815.835 -4.245 816.165 -3.915 ;
        RECT 814.475 -4.245 814.805 -3.915 ;
        RECT 813.115 -4.245 813.445 -3.915 ;
        RECT 811.755 -4.245 812.085 -3.915 ;
        RECT 810.395 -4.245 810.725 -3.915 ;
        RECT 809.035 -4.245 809.365 -3.915 ;
        RECT 807.675 -4.245 808.005 -3.915 ;
        RECT 806.315 -4.245 806.645 -3.915 ;
        RECT 804.955 -4.245 805.285 -3.915 ;
        RECT 803.595 -4.245 803.925 -3.915 ;
        RECT 802.235 -4.245 802.565 -3.915 ;
        RECT 800.875 -4.245 801.205 -3.915 ;
        RECT 799.515 -4.245 799.845 -3.915 ;
        RECT 798.155 -4.245 798.485 -3.915 ;
        RECT 796.795 -4.245 797.125 -3.915 ;
        RECT 795.435 -4.245 795.765 -3.915 ;
        RECT 794.075 -4.245 794.405 -3.915 ;
        RECT 792.715 -4.245 793.045 -3.915 ;
        RECT 791.355 -4.245 791.685 -3.915 ;
        RECT 789.995 -4.245 790.325 -3.915 ;
        RECT 788.635 -4.245 788.965 -3.915 ;
        RECT 787.275 -4.245 787.605 -3.915 ;
        RECT 785.915 -4.245 786.245 -3.915 ;
        RECT 784.555 -4.245 784.885 -3.915 ;
        RECT 783.195 -4.245 783.525 -3.915 ;
        RECT 781.835 -4.245 782.165 -3.915 ;
        RECT 780.475 -4.245 780.805 -3.915 ;
        RECT 779.115 -4.245 779.445 -3.915 ;
        RECT 777.755 -4.245 778.085 -3.915 ;
        RECT 776.395 -4.245 776.725 -3.915 ;
        RECT 775.035 -4.245 775.365 -3.915 ;
        RECT 773.675 -4.245 774.005 -3.915 ;
        RECT 772.315 -4.245 772.645 -3.915 ;
        RECT 770.955 -4.245 771.285 -3.915 ;
        RECT 769.595 -4.245 769.925 -3.915 ;
        RECT 768.235 -4.245 768.565 -3.915 ;
        RECT 766.875 -4.245 767.205 -3.915 ;
        RECT 765.515 -4.245 765.845 -3.915 ;
        RECT 764.155 -4.245 764.485 -3.915 ;
        RECT 762.795 -4.245 763.125 -3.915 ;
        RECT 761.435 -4.245 761.765 -3.915 ;
        RECT 760.075 -4.245 760.405 -3.915 ;
        RECT 758.715 -4.245 759.045 -3.915 ;
        RECT 757.355 -4.245 757.685 -3.915 ;
        RECT 755.995 -4.245 756.325 -3.915 ;
        RECT 754.635 -4.245 754.965 -3.915 ;
        RECT 753.275 -4.245 753.605 -3.915 ;
        RECT 751.915 -4.245 752.245 -3.915 ;
        RECT 750.555 -4.245 750.885 -3.915 ;
        RECT 749.195 -4.245 749.525 -3.915 ;
        RECT 747.835 -4.245 748.165 -3.915 ;
        RECT 746.475 -4.245 746.805 -3.915 ;
        RECT 745.115 -4.245 745.445 -3.915 ;
        RECT 743.755 -4.245 744.085 -3.915 ;
        RECT 742.395 -4.245 742.725 -3.915 ;
        RECT 741.035 -4.245 741.365 -3.915 ;
        RECT 739.675 -4.245 740.005 -3.915 ;
        RECT 738.315 -4.245 738.645 -3.915 ;
        RECT 736.955 -4.245 737.285 -3.915 ;
        RECT 735.595 -4.245 735.925 -3.915 ;
        RECT 734.235 -4.245 734.565 -3.915 ;
        RECT 732.875 -4.245 733.205 -3.915 ;
        RECT 731.515 -4.245 731.845 -3.915 ;
        RECT 730.155 -4.245 730.485 -3.915 ;
        RECT 728.795 -4.245 729.125 -3.915 ;
        RECT 727.435 -4.245 727.765 -3.915 ;
        RECT 726.075 -4.245 726.405 -3.915 ;
        RECT 724.715 -4.245 725.045 -3.915 ;
        RECT 723.355 -4.245 723.685 -3.915 ;
        RECT 721.995 -4.245 722.325 -3.915 ;
        RECT 720.635 -4.245 720.965 -3.915 ;
        RECT 719.275 -4.245 719.605 -3.915 ;
        RECT 717.915 -4.245 718.245 -3.915 ;
        RECT 716.555 -4.245 716.885 -3.915 ;
        RECT 715.195 -4.245 715.525 -3.915 ;
        RECT 713.835 -4.245 714.165 -3.915 ;
        RECT 712.475 -4.245 712.805 -3.915 ;
        RECT 711.115 -4.245 711.445 -3.915 ;
        RECT 709.755 -4.245 710.085 -3.915 ;
        RECT 708.395 -4.245 708.725 -3.915 ;
        RECT 707.035 -4.245 707.365 -3.915 ;
        RECT 705.675 -4.245 706.005 -3.915 ;
        RECT 704.315 -4.245 704.645 -3.915 ;
        RECT 702.955 -4.245 703.285 -3.915 ;
        RECT 701.595 -4.245 701.925 -3.915 ;
        RECT 700.235 -4.245 700.565 -3.915 ;
        RECT 698.875 -4.245 699.205 -3.915 ;
        RECT 697.515 -4.245 697.845 -3.915 ;
        RECT 696.155 -4.245 696.485 -3.915 ;
        RECT 694.795 -4.245 695.125 -3.915 ;
        RECT 693.435 -4.245 693.765 -3.915 ;
        RECT 692.075 -4.245 692.405 -3.915 ;
        RECT 690.715 -4.245 691.045 -3.915 ;
        RECT 689.355 -4.245 689.685 -3.915 ;
        RECT 687.995 -4.245 688.325 -3.915 ;
        RECT 686.635 -4.245 686.965 -3.915 ;
        RECT 685.275 -4.245 685.605 -3.915 ;
        RECT 683.915 -4.245 684.245 -3.915 ;
        RECT 682.555 -4.245 682.885 -3.915 ;
        RECT 681.195 -4.245 681.525 -3.915 ;
        RECT 679.835 -4.245 680.165 -3.915 ;
        RECT 678.475 -4.245 678.805 -3.915 ;
        RECT 954.555 -4.245 954.885 -3.915 ;
        RECT 678.475 -4.24 954.885 -3.92 ;
        RECT 953.195 -4.245 953.525 -3.915 ;
        RECT 951.835 -4.245 952.165 -3.915 ;
        RECT 950.475 -4.245 950.805 -3.915 ;
        RECT 949.115 -4.245 949.445 -3.915 ;
        RECT 947.755 -4.245 948.085 -3.915 ;
        RECT 946.395 -4.245 946.725 -3.915 ;
        RECT 945.035 -4.245 945.365 -3.915 ;
        RECT 943.675 -4.245 944.005 -3.915 ;
        RECT 942.315 -4.245 942.645 -3.915 ;
        RECT 940.955 -4.245 941.285 -3.915 ;
        RECT 939.595 -4.245 939.925 -3.915 ;
        RECT 938.235 -4.245 938.565 -3.915 ;
        RECT 936.875 -4.245 937.205 -3.915 ;
        RECT 935.515 -4.245 935.845 -3.915 ;
        RECT 934.155 -4.245 934.485 -3.915 ;
        RECT 932.795 -4.245 933.125 -3.915 ;
        RECT 931.435 -4.245 931.765 -3.915 ;
        RECT 930.075 -4.245 930.405 -3.915 ;
        RECT 928.715 -4.245 929.045 -3.915 ;
        RECT 927.355 -4.245 927.685 -3.915 ;
        RECT 925.995 -4.245 926.325 -3.915 ;
        RECT 924.635 -4.245 924.965 -3.915 ;
        RECT 923.275 -4.245 923.605 -3.915 ;
        RECT 921.915 -4.245 922.245 -3.915 ;
        RECT 920.555 -4.245 920.885 -3.915 ;
        RECT 919.195 -4.245 919.525 -3.915 ;
        RECT 917.835 -4.245 918.165 -3.915 ;
        RECT 916.475 -4.245 916.805 -3.915 ;
        RECT 915.115 -4.245 915.445 -3.915 ;
        RECT 913.755 -4.245 914.085 -3.915 ;
        RECT 912.395 -4.245 912.725 -3.915 ;
        RECT 911.035 -4.245 911.365 -3.915 ;
        RECT 909.675 -4.245 910.005 -3.915 ;
        RECT 908.315 -4.245 908.645 -3.915 ;
        RECT 906.955 -4.245 907.285 -3.915 ;
        RECT 905.595 -4.245 905.925 -3.915 ;
        RECT 904.235 -4.245 904.565 -3.915 ;
        RECT 902.875 -4.245 903.205 -3.915 ;
        RECT 901.515 -4.245 901.845 -3.915 ;
        RECT 900.155 -4.245 900.485 -3.915 ;
        RECT 898.795 -4.245 899.125 -3.915 ;
        RECT 897.435 -4.245 897.765 -3.915 ;
        RECT 896.075 -4.245 896.405 -3.915 ;
        RECT 894.715 -4.245 895.045 -3.915 ;
        RECT 893.355 -4.245 893.685 -3.915 ;
        RECT 891.995 -4.245 892.325 -3.915 ;
        RECT 890.635 -4.245 890.965 -3.915 ;
        RECT 889.275 -4.245 889.605 -3.915 ;
        RECT 887.915 -4.245 888.245 -3.915 ;
        RECT 886.555 -4.245 886.885 -3.915 ;
        RECT 885.195 -4.245 885.525 -3.915 ;
        RECT 883.835 -4.245 884.165 -3.915 ;
        RECT 882.475 -4.245 882.805 -3.915 ;
        RECT 881.115 -4.245 881.445 -3.915 ;
        RECT 879.755 -4.245 880.085 -3.915 ;
        RECT 878.395 -4.245 878.725 -3.915 ;
        RECT 877.035 -4.245 877.365 -3.915 ;
        RECT 875.675 -4.245 876.005 -3.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 653.995 -5.605 654.325 -5.275 ;
        RECT 652.635 -5.605 652.965 -5.275 ;
        RECT 651.275 -5.605 651.605 -5.275 ;
        RECT 649.915 -5.605 650.245 -5.275 ;
        RECT 648.555 -5.605 648.885 -5.275 ;
        RECT 647.195 -5.605 647.525 -5.275 ;
        RECT 645.835 -5.605 646.165 -5.275 ;
        RECT 644.475 -5.605 644.805 -5.275 ;
        RECT 643.115 -5.605 643.445 -5.275 ;
        RECT 641.755 -5.605 642.085 -5.275 ;
        RECT 640.395 -5.605 640.725 -5.275 ;
        RECT 639.035 -5.605 639.365 -5.275 ;
        RECT 637.675 -5.605 638.005 -5.275 ;
        RECT 636.315 -5.605 636.645 -5.275 ;
        RECT 634.955 -5.605 635.285 -5.275 ;
        RECT 633.595 -5.605 633.925 -5.275 ;
        RECT 632.235 -5.605 632.565 -5.275 ;
        RECT 630.875 -5.605 631.205 -5.275 ;
        RECT 629.515 -5.605 629.845 -5.275 ;
        RECT 628.155 -5.605 628.485 -5.275 ;
        RECT 626.795 -5.605 627.125 -5.275 ;
        RECT 625.435 -5.605 625.765 -5.275 ;
        RECT 624.075 -5.605 624.405 -5.275 ;
        RECT 622.715 -5.605 623.045 -5.275 ;
        RECT 621.355 -5.605 621.685 -5.275 ;
        RECT 619.995 -5.605 620.325 -5.275 ;
        RECT 618.635 -5.605 618.965 -5.275 ;
        RECT 617.275 -5.605 617.605 -5.275 ;
        RECT 615.915 -5.605 616.245 -5.275 ;
        RECT 614.555 -5.605 614.885 -5.275 ;
        RECT 613.195 -5.605 613.525 -5.275 ;
        RECT 611.835 -5.605 612.165 -5.275 ;
        RECT 610.475 -5.605 610.805 -5.275 ;
        RECT 609.115 -5.605 609.445 -5.275 ;
        RECT 607.755 -5.605 608.085 -5.275 ;
        RECT 606.395 -5.605 606.725 -5.275 ;
        RECT 605.035 -5.605 605.365 -5.275 ;
        RECT 603.675 -5.605 604.005 -5.275 ;
        RECT 602.315 -5.605 602.645 -5.275 ;
        RECT 600.955 -5.605 601.285 -5.275 ;
        RECT 599.595 -5.605 599.925 -5.275 ;
        RECT 598.235 -5.605 598.565 -5.275 ;
        RECT 596.875 -5.605 597.205 -5.275 ;
        RECT 595.515 -5.605 595.845 -5.275 ;
        RECT 594.155 -5.605 594.485 -5.275 ;
        RECT 592.795 -5.605 593.125 -5.275 ;
        RECT 591.435 -5.605 591.765 -5.275 ;
        RECT 590.075 -5.605 590.405 -5.275 ;
        RECT 588.715 -5.605 589.045 -5.275 ;
        RECT 587.355 -5.605 587.685 -5.275 ;
        RECT 585.995 -5.605 586.325 -5.275 ;
        RECT 584.635 -5.605 584.965 -5.275 ;
        RECT 583.275 -5.605 583.605 -5.275 ;
        RECT 581.915 -5.605 582.245 -5.275 ;
        RECT 580.555 -5.605 580.885 -5.275 ;
        RECT 579.195 -5.605 579.525 -5.275 ;
        RECT 577.835 -5.605 578.165 -5.275 ;
        RECT 576.475 -5.605 576.805 -5.275 ;
        RECT 575.115 -5.605 575.445 -5.275 ;
        RECT 573.755 -5.605 574.085 -5.275 ;
        RECT 572.395 -5.605 572.725 -5.275 ;
        RECT 571.035 -5.605 571.365 -5.275 ;
        RECT 569.675 -5.605 570.005 -5.275 ;
        RECT 568.315 -5.605 568.645 -5.275 ;
        RECT 566.955 -5.605 567.285 -5.275 ;
        RECT 565.595 -5.605 565.925 -5.275 ;
        RECT 564.235 -5.605 564.565 -5.275 ;
        RECT 562.875 -5.605 563.205 -5.275 ;
        RECT 561.515 -5.605 561.845 -5.275 ;
        RECT 560.155 -5.605 560.485 -5.275 ;
        RECT 558.795 -5.605 559.125 -5.275 ;
        RECT 557.435 -5.605 557.765 -5.275 ;
        RECT 556.075 -5.605 556.405 -5.275 ;
        RECT 554.715 -5.605 555.045 -5.275 ;
        RECT 553.355 -5.605 553.685 -5.275 ;
        RECT 551.995 -5.605 552.325 -5.275 ;
        RECT 550.635 -5.605 550.965 -5.275 ;
        RECT 549.275 -5.605 549.605 -5.275 ;
        RECT 547.915 -5.605 548.245 -5.275 ;
        RECT 546.555 -5.605 546.885 -5.275 ;
        RECT 545.195 -5.605 545.525 -5.275 ;
        RECT 543.835 -5.605 544.165 -5.275 ;
        RECT 542.475 -5.605 542.805 -5.275 ;
        RECT 541.115 -5.605 541.445 -5.275 ;
        RECT 539.755 -5.605 540.085 -5.275 ;
        RECT 538.395 -5.605 538.725 -5.275 ;
        RECT 537.035 -5.605 537.365 -5.275 ;
        RECT 535.675 -5.605 536.005 -5.275 ;
        RECT 534.315 -5.605 534.645 -5.275 ;
        RECT 532.955 -5.605 533.285 -5.275 ;
        RECT 531.595 -5.605 531.925 -5.275 ;
        RECT 530.235 -5.605 530.565 -5.275 ;
        RECT 528.875 -5.605 529.205 -5.275 ;
        RECT 527.515 -5.605 527.845 -5.275 ;
        RECT 526.155 -5.605 526.485 -5.275 ;
        RECT 524.795 -5.605 525.125 -5.275 ;
        RECT 523.435 -5.605 523.765 -5.275 ;
        RECT 522.075 -5.605 522.405 -5.275 ;
        RECT 520.715 -5.605 521.045 -5.275 ;
        RECT 519.355 -5.605 519.685 -5.275 ;
        RECT 517.995 -5.605 518.325 -5.275 ;
        RECT 516.635 -5.605 516.965 -5.275 ;
        RECT 515.275 -5.605 515.605 -5.275 ;
        RECT 513.915 -5.605 514.245 -5.275 ;
        RECT 512.555 -5.605 512.885 -5.275 ;
        RECT 511.195 -5.605 511.525 -5.275 ;
        RECT 509.835 -5.605 510.165 -5.275 ;
        RECT 508.475 -5.605 508.805 -5.275 ;
        RECT 507.115 -5.605 507.445 -5.275 ;
        RECT 505.755 -5.605 506.085 -5.275 ;
        RECT 504.395 -5.605 504.725 -5.275 ;
        RECT 503.035 -5.605 503.365 -5.275 ;
        RECT 501.675 -5.605 502.005 -5.275 ;
        RECT 500.315 -5.605 500.645 -5.275 ;
        RECT 498.955 -5.605 499.285 -5.275 ;
        RECT 497.595 -5.605 497.925 -5.275 ;
        RECT 496.235 -5.605 496.565 -5.275 ;
        RECT 494.875 -5.605 495.205 -5.275 ;
        RECT 493.515 -5.605 493.845 -5.275 ;
        RECT 492.155 -5.605 492.485 -5.275 ;
        RECT 490.795 -5.605 491.125 -5.275 ;
        RECT 489.435 -5.605 489.765 -5.275 ;
        RECT 488.075 -5.605 488.405 -5.275 ;
        RECT 486.715 -5.605 487.045 -5.275 ;
        RECT 485.355 -5.605 485.685 -5.275 ;
        RECT 483.995 -5.605 484.325 -5.275 ;
        RECT 482.635 -5.605 482.965 -5.275 ;
        RECT 481.275 -5.605 481.605 -5.275 ;
        RECT 479.915 -5.605 480.245 -5.275 ;
        RECT 478.555 -5.605 478.885 -5.275 ;
        RECT 477.195 -5.605 477.525 -5.275 ;
        RECT 475.835 -5.605 476.165 -5.275 ;
        RECT 474.475 -5.605 474.805 -5.275 ;
        RECT 473.115 -5.605 473.445 -5.275 ;
        RECT 471.755 -5.605 472.085 -5.275 ;
        RECT 470.395 -5.605 470.725 -5.275 ;
        RECT 469.035 -5.605 469.365 -5.275 ;
        RECT 467.675 -5.605 468.005 -5.275 ;
        RECT 466.315 -5.605 466.645 -5.275 ;
        RECT 464.955 -5.605 465.285 -5.275 ;
        RECT 463.595 -5.605 463.925 -5.275 ;
        RECT 462.235 -5.605 462.565 -5.275 ;
        RECT 460.875 -5.605 461.205 -5.275 ;
        RECT 459.515 -5.605 459.845 -5.275 ;
        RECT 458.155 -5.605 458.485 -5.275 ;
        RECT 456.795 -5.605 457.125 -5.275 ;
        RECT 455.435 -5.605 455.765 -5.275 ;
        RECT 454.075 -5.605 454.405 -5.275 ;
        RECT 452.715 -5.605 453.045 -5.275 ;
        RECT 451.355 -5.605 451.685 -5.275 ;
        RECT 449.995 -5.605 450.325 -5.275 ;
        RECT 448.635 -5.605 448.965 -5.275 ;
        RECT 447.275 -5.605 447.605 -5.275 ;
        RECT 445.915 -5.605 446.245 -5.275 ;
        RECT 444.555 -5.605 444.885 -5.275 ;
        RECT 443.195 -5.605 443.525 -5.275 ;
        RECT 441.835 -5.605 442.165 -5.275 ;
        RECT 440.475 -5.605 440.805 -5.275 ;
        RECT 439.115 -5.605 439.445 -5.275 ;
        RECT 437.755 -5.605 438.085 -5.275 ;
        RECT 436.395 -5.605 436.725 -5.275 ;
        RECT 435.035 -5.605 435.365 -5.275 ;
        RECT 433.675 -5.605 434.005 -5.275 ;
        RECT 432.315 -5.605 432.645 -5.275 ;
        RECT 430.955 -5.605 431.285 -5.275 ;
        RECT 429.595 -5.605 429.925 -5.275 ;
        RECT 428.235 -5.605 428.565 -5.275 ;
        RECT 426.875 -5.605 427.205 -5.275 ;
        RECT 425.515 -5.605 425.845 -5.275 ;
        RECT 424.155 -5.605 424.485 -5.275 ;
        RECT 422.795 -5.605 423.125 -5.275 ;
        RECT 421.435 -5.605 421.765 -5.275 ;
        RECT 420.075 -5.605 420.405 -5.275 ;
        RECT 418.715 -5.605 419.045 -5.275 ;
        RECT 417.355 -5.605 417.685 -5.275 ;
        RECT 415.995 -5.605 416.325 -5.275 ;
        RECT 414.635 -5.605 414.965 -5.275 ;
        RECT 413.275 -5.605 413.605 -5.275 ;
        RECT 411.915 -5.605 412.245 -5.275 ;
        RECT 410.555 -5.605 410.885 -5.275 ;
        RECT 409.195 -5.605 409.525 -5.275 ;
        RECT 407.835 -5.605 408.165 -5.275 ;
        RECT 406.475 -5.605 406.805 -5.275 ;
        RECT 405.115 -5.605 405.445 -5.275 ;
        RECT 403.755 -5.605 404.085 -5.275 ;
        RECT 402.395 -5.605 402.725 -5.275 ;
        RECT 401.035 -5.605 401.365 -5.275 ;
        RECT 399.675 -5.605 400.005 -5.275 ;
        RECT 398.315 -5.605 398.645 -5.275 ;
        RECT 396.955 -5.605 397.285 -5.275 ;
        RECT 395.595 -5.605 395.925 -5.275 ;
        RECT 394.235 -5.605 394.565 -5.275 ;
        RECT 392.875 -5.605 393.205 -5.275 ;
        RECT 391.515 -5.605 391.845 -5.275 ;
        RECT 390.155 -5.605 390.485 -5.275 ;
        RECT 388.795 -5.605 389.125 -5.275 ;
        RECT 387.435 -5.605 387.765 -5.275 ;
        RECT 386.075 -5.605 386.405 -5.275 ;
        RECT 384.715 -5.605 385.045 -5.275 ;
        RECT 383.355 -5.605 383.685 -5.275 ;
        RECT 381.995 -5.605 382.325 -5.275 ;
        RECT 380.635 -5.605 380.965 -5.275 ;
        RECT 379.275 -5.605 379.605 -5.275 ;
        RECT 377.915 -5.605 378.245 -5.275 ;
        RECT 376.555 -5.605 376.885 -5.275 ;
        RECT 375.195 -5.605 375.525 -5.275 ;
        RECT 373.835 -5.605 374.165 -5.275 ;
        RECT 372.475 -5.605 372.805 -5.275 ;
        RECT 371.115 -5.605 371.445 -5.275 ;
        RECT 369.755 -5.605 370.085 -5.275 ;
        RECT 368.395 -5.605 368.725 -5.275 ;
        RECT 367.035 -5.605 367.365 -5.275 ;
        RECT 365.675 -5.605 366.005 -5.275 ;
        RECT 364.315 -5.605 364.645 -5.275 ;
        RECT 362.955 -5.605 363.285 -5.275 ;
        RECT 361.595 -5.605 361.925 -5.275 ;
        RECT 360.235 -5.605 360.565 -5.275 ;
        RECT 358.875 -5.605 359.205 -5.275 ;
        RECT 357.515 -5.605 357.845 -5.275 ;
        RECT 356.155 -5.605 356.485 -5.275 ;
        RECT 354.795 -5.605 355.125 -5.275 ;
        RECT 353.435 -5.605 353.765 -5.275 ;
        RECT 352.075 -5.605 352.405 -5.275 ;
        RECT 350.715 -5.605 351.045 -5.275 ;
        RECT 349.355 -5.605 349.685 -5.275 ;
        RECT 347.995 -5.605 348.325 -5.275 ;
        RECT 346.635 -5.605 346.965 -5.275 ;
        RECT 345.275 -5.605 345.605 -5.275 ;
        RECT 343.915 -5.605 344.245 -5.275 ;
        RECT 342.555 -5.605 342.885 -5.275 ;
        RECT 341.195 -5.605 341.525 -5.275 ;
        RECT 339.835 -5.605 340.165 -5.275 ;
        RECT 338.475 -5.605 338.805 -5.275 ;
        RECT 337.115 -5.605 337.445 -5.275 ;
        RECT 335.755 -5.605 336.085 -5.275 ;
        RECT 334.395 -5.605 334.725 -5.275 ;
        RECT 333.035 -5.605 333.365 -5.275 ;
        RECT 331.675 -5.605 332.005 -5.275 ;
        RECT 330.315 -5.605 330.645 -5.275 ;
        RECT 328.955 -5.605 329.285 -5.275 ;
        RECT 327.595 -5.605 327.925 -5.275 ;
        RECT 326.235 -5.605 326.565 -5.275 ;
        RECT 324.875 -5.605 325.205 -5.275 ;
        RECT 323.515 -5.605 323.845 -5.275 ;
        RECT 322.155 -5.605 322.485 -5.275 ;
        RECT 320.795 -5.605 321.125 -5.275 ;
        RECT 319.435 -5.605 319.765 -5.275 ;
        RECT 318.075 -5.605 318.405 -5.275 ;
        RECT 316.715 -5.605 317.045 -5.275 ;
        RECT 315.355 -5.605 315.685 -5.275 ;
        RECT 313.995 -5.605 314.325 -5.275 ;
        RECT 312.635 -5.605 312.965 -5.275 ;
        RECT 311.275 -5.605 311.605 -5.275 ;
        RECT 309.915 -5.605 310.245 -5.275 ;
        RECT 308.555 -5.605 308.885 -5.275 ;
        RECT 307.195 -5.605 307.525 -5.275 ;
        RECT 305.835 -5.605 306.165 -5.275 ;
        RECT 304.475 -5.605 304.805 -5.275 ;
        RECT 303.115 -5.605 303.445 -5.275 ;
        RECT 301.755 -5.605 302.085 -5.275 ;
        RECT 300.395 -5.605 300.725 -5.275 ;
        RECT 299.035 -5.605 299.365 -5.275 ;
        RECT 297.675 -5.605 298.005 -5.275 ;
        RECT 296.315 -5.605 296.645 -5.275 ;
        RECT 294.955 -5.605 295.285 -5.275 ;
        RECT 293.595 -5.605 293.925 -5.275 ;
        RECT 292.235 -5.605 292.565 -5.275 ;
        RECT 290.875 -5.605 291.205 -5.275 ;
        RECT 289.515 -5.605 289.845 -5.275 ;
        RECT 288.155 -5.605 288.485 -5.275 ;
        RECT 286.795 -5.605 287.125 -5.275 ;
        RECT 285.435 -5.605 285.765 -5.275 ;
        RECT 284.075 -5.605 284.405 -5.275 ;
        RECT 282.715 -5.605 283.045 -5.275 ;
        RECT 281.355 -5.605 281.685 -5.275 ;
        RECT 279.995 -5.605 280.325 -5.275 ;
        RECT 278.635 -5.605 278.965 -5.275 ;
        RECT 277.275 -5.605 277.605 -5.275 ;
        RECT 275.915 -5.605 276.245 -5.275 ;
        RECT 274.555 -5.605 274.885 -5.275 ;
        RECT 273.195 -5.605 273.525 -5.275 ;
        RECT 271.835 -5.605 272.165 -5.275 ;
        RECT 270.475 -5.605 270.805 -5.275 ;
        RECT 269.115 -5.605 269.445 -5.275 ;
        RECT 267.755 -5.605 268.085 -5.275 ;
        RECT 266.395 -5.605 266.725 -5.275 ;
        RECT 265.035 -5.605 265.365 -5.275 ;
        RECT 263.675 -5.605 264.005 -5.275 ;
        RECT 262.315 -5.605 262.645 -5.275 ;
        RECT 260.955 -5.605 261.285 -5.275 ;
        RECT 259.595 -5.605 259.925 -5.275 ;
        RECT 258.235 -5.605 258.565 -5.275 ;
        RECT 256.875 -5.605 257.205 -5.275 ;
        RECT 255.515 -5.605 255.845 -5.275 ;
        RECT 254.155 -5.605 254.485 -5.275 ;
        RECT 252.795 -5.605 253.125 -5.275 ;
        RECT 251.435 -5.605 251.765 -5.275 ;
        RECT 250.075 -5.605 250.405 -5.275 ;
        RECT 248.715 -5.605 249.045 -5.275 ;
        RECT 247.355 -5.605 247.685 -5.275 ;
        RECT 245.995 -5.605 246.325 -5.275 ;
        RECT 244.635 -5.605 244.965 -5.275 ;
        RECT 243.275 -5.605 243.605 -5.275 ;
        RECT 241.915 -5.605 242.245 -5.275 ;
        RECT 240.555 -5.605 240.885 -5.275 ;
        RECT 239.195 -5.605 239.525 -5.275 ;
        RECT 237.835 -5.605 238.165 -5.275 ;
        RECT 236.475 -5.605 236.805 -5.275 ;
        RECT 235.115 -5.605 235.445 -5.275 ;
        RECT 233.755 -5.605 234.085 -5.275 ;
        RECT 232.395 -5.605 232.725 -5.275 ;
        RECT 231.035 -5.605 231.365 -5.275 ;
        RECT 229.675 -5.605 230.005 -5.275 ;
        RECT 228.315 -5.605 228.645 -5.275 ;
        RECT 226.955 -5.605 227.285 -5.275 ;
        RECT 225.595 -5.605 225.925 -5.275 ;
        RECT 224.235 -5.605 224.565 -5.275 ;
        RECT 222.875 -5.605 223.205 -5.275 ;
        RECT 221.515 -5.605 221.845 -5.275 ;
        RECT 220.155 -5.605 220.485 -5.275 ;
        RECT 218.795 -5.605 219.125 -5.275 ;
        RECT 217.435 -5.605 217.765 -5.275 ;
        RECT 216.075 -5.605 216.405 -5.275 ;
        RECT 214.715 -5.605 215.045 -5.275 ;
        RECT 213.355 -5.605 213.685 -5.275 ;
        RECT 211.995 -5.605 212.325 -5.275 ;
        RECT 210.635 -5.605 210.965 -5.275 ;
        RECT 209.275 -5.605 209.605 -5.275 ;
        RECT 207.915 -5.605 208.245 -5.275 ;
        RECT 206.555 -5.605 206.885 -5.275 ;
        RECT 205.195 -5.605 205.525 -5.275 ;
        RECT 203.835 -5.605 204.165 -5.275 ;
        RECT 202.475 -5.605 202.805 -5.275 ;
        RECT 201.115 -5.605 201.445 -5.275 ;
        RECT 199.755 -5.605 200.085 -5.275 ;
        RECT 198.395 -5.605 198.725 -5.275 ;
        RECT 197.035 -5.605 197.365 -5.275 ;
        RECT 195.675 -5.605 196.005 -5.275 ;
        RECT 194.315 -5.605 194.645 -5.275 ;
        RECT 192.955 -5.605 193.285 -5.275 ;
        RECT 191.595 -5.605 191.925 -5.275 ;
        RECT 190.235 -5.605 190.565 -5.275 ;
        RECT 188.875 -5.605 189.205 -5.275 ;
        RECT 187.515 -5.605 187.845 -5.275 ;
        RECT 186.155 -5.605 186.485 -5.275 ;
        RECT 184.795 -5.605 185.125 -5.275 ;
        RECT 183.435 -5.605 183.765 -5.275 ;
        RECT 182.075 -5.605 182.405 -5.275 ;
        RECT 180.715 -5.605 181.045 -5.275 ;
        RECT 179.355 -5.605 179.685 -5.275 ;
        RECT 177.995 -5.605 178.325 -5.275 ;
        RECT 176.635 -5.605 176.965 -5.275 ;
        RECT 175.275 -5.605 175.605 -5.275 ;
        RECT 173.915 -5.605 174.245 -5.275 ;
        RECT 172.555 -5.605 172.885 -5.275 ;
        RECT 171.195 -5.605 171.525 -5.275 ;
        RECT 169.835 -5.605 170.165 -5.275 ;
        RECT 168.475 -5.605 168.805 -5.275 ;
        RECT 167.115 -5.605 167.445 -5.275 ;
        RECT 165.755 -5.605 166.085 -5.275 ;
        RECT 164.395 -5.605 164.725 -5.275 ;
        RECT 163.035 -5.605 163.365 -5.275 ;
        RECT 161.675 -5.605 162.005 -5.275 ;
        RECT 160.315 -5.605 160.645 -5.275 ;
        RECT 158.955 -5.605 159.285 -5.275 ;
        RECT 157.595 -5.605 157.925 -5.275 ;
        RECT 156.235 -5.605 156.565 -5.275 ;
        RECT 154.875 -5.605 155.205 -5.275 ;
        RECT 153.515 -5.605 153.845 -5.275 ;
        RECT 152.155 -5.605 152.485 -5.275 ;
        RECT 150.795 -5.605 151.125 -5.275 ;
        RECT 149.435 -5.605 149.765 -5.275 ;
        RECT 148.075 -5.605 148.405 -5.275 ;
        RECT 146.715 -5.605 147.045 -5.275 ;
        RECT 145.355 -5.605 145.685 -5.275 ;
        RECT 143.995 -5.605 144.325 -5.275 ;
        RECT 142.635 -5.605 142.965 -5.275 ;
        RECT 141.275 -5.605 141.605 -5.275 ;
        RECT 139.915 -5.605 140.245 -5.275 ;
        RECT 138.555 -5.605 138.885 -5.275 ;
        RECT 137.195 -5.605 137.525 -5.275 ;
        RECT 135.835 -5.605 136.165 -5.275 ;
        RECT 134.475 -5.605 134.805 -5.275 ;
        RECT 133.115 -5.605 133.445 -5.275 ;
        RECT 131.755 -5.605 132.085 -5.275 ;
        RECT 130.395 -5.605 130.725 -5.275 ;
        RECT 129.035 -5.605 129.365 -5.275 ;
        RECT 127.675 -5.605 128.005 -5.275 ;
        RECT 126.315 -5.605 126.645 -5.275 ;
        RECT 124.955 -5.605 125.285 -5.275 ;
        RECT 123.595 -5.605 123.925 -5.275 ;
        RECT 122.235 -5.605 122.565 -5.275 ;
        RECT 120.875 -5.605 121.205 -5.275 ;
        RECT 119.515 -5.605 119.845 -5.275 ;
        RECT 118.155 -5.605 118.485 -5.275 ;
        RECT 116.795 -5.605 117.125 -5.275 ;
        RECT 115.435 -5.605 115.765 -5.275 ;
        RECT 114.075 -5.605 114.405 -5.275 ;
        RECT 112.715 -5.605 113.045 -5.275 ;
        RECT 111.355 -5.605 111.685 -5.275 ;
        RECT 109.995 -5.605 110.325 -5.275 ;
        RECT 108.635 -5.605 108.965 -5.275 ;
        RECT 107.275 -5.605 107.605 -5.275 ;
        RECT 105.915 -5.605 106.245 -5.275 ;
        RECT 104.555 -5.605 104.885 -5.275 ;
        RECT 103.195 -5.605 103.525 -5.275 ;
        RECT 101.835 -5.605 102.165 -5.275 ;
        RECT 100.475 -5.605 100.805 -5.275 ;
        RECT 99.115 -5.605 99.445 -5.275 ;
        RECT 97.755 -5.605 98.085 -5.275 ;
        RECT 96.395 -5.605 96.725 -5.275 ;
        RECT 95.035 -5.605 95.365 -5.275 ;
        RECT 93.675 -5.605 94.005 -5.275 ;
        RECT 92.315 -5.605 92.645 -5.275 ;
        RECT 90.955 -5.605 91.285 -5.275 ;
        RECT 89.595 -5.605 89.925 -5.275 ;
        RECT 88.235 -5.605 88.565 -5.275 ;
        RECT 86.875 -5.605 87.205 -5.275 ;
        RECT 85.515 -5.605 85.845 -5.275 ;
        RECT 84.155 -5.605 84.485 -5.275 ;
        RECT 82.795 -5.605 83.125 -5.275 ;
        RECT 81.435 -5.605 81.765 -5.275 ;
        RECT 80.075 -5.605 80.405 -5.275 ;
        RECT 78.715 -5.605 79.045 -5.275 ;
        RECT 77.355 -5.605 77.685 -5.275 ;
        RECT 75.995 -5.605 76.325 -5.275 ;
        RECT 74.635 -5.605 74.965 -5.275 ;
        RECT 73.275 -5.605 73.605 -5.275 ;
        RECT 71.915 -5.605 72.245 -5.275 ;
        RECT 70.555 -5.605 70.885 -5.275 ;
        RECT 69.195 -5.605 69.525 -5.275 ;
        RECT 67.835 -5.605 68.165 -5.275 ;
        RECT 66.475 -5.605 66.805 -5.275 ;
        RECT 65.115 -5.605 65.445 -5.275 ;
        RECT 63.755 -5.605 64.085 -5.275 ;
        RECT 62.395 -5.605 62.725 -5.275 ;
        RECT 61.035 -5.605 61.365 -5.275 ;
        RECT 59.675 -5.605 60.005 -5.275 ;
        RECT 58.315 -5.605 58.645 -5.275 ;
        RECT 56.955 -5.605 57.285 -5.275 ;
        RECT 55.595 -5.605 55.925 -5.275 ;
        RECT 54.235 -5.605 54.565 -5.275 ;
        RECT 52.875 -5.605 53.205 -5.275 ;
        RECT 51.515 -5.605 51.845 -5.275 ;
        RECT 50.155 -5.605 50.485 -5.275 ;
        RECT 48.795 -5.605 49.125 -5.275 ;
        RECT 47.435 -5.605 47.765 -5.275 ;
        RECT 46.075 -5.605 46.405 -5.275 ;
        RECT 44.715 -5.605 45.045 -5.275 ;
        RECT 43.355 -5.605 43.685 -5.275 ;
        RECT 41.995 -5.605 42.325 -5.275 ;
        RECT 40.635 -5.605 40.965 -5.275 ;
        RECT 39.275 -5.605 39.605 -5.275 ;
        RECT 37.915 -5.605 38.245 -5.275 ;
        RECT 36.555 -5.605 36.885 -5.275 ;
        RECT 35.195 -5.605 35.525 -5.275 ;
        RECT 33.835 -5.605 34.165 -5.275 ;
        RECT 32.475 -5.605 32.805 -5.275 ;
        RECT 31.115 -5.605 31.445 -5.275 ;
        RECT 29.755 -5.605 30.085 -5.275 ;
        RECT 28.395 -5.605 28.725 -5.275 ;
        RECT 27.035 -5.605 27.365 -5.275 ;
        RECT 25.675 -5.605 26.005 -5.275 ;
        RECT 24.315 -5.605 24.645 -5.275 ;
        RECT 22.955 -5.605 23.285 -5.275 ;
        RECT 21.595 -5.605 21.925 -5.275 ;
        RECT 20.235 -5.605 20.565 -5.275 ;
        RECT 18.875 -5.605 19.205 -5.275 ;
        RECT 17.515 -5.605 17.845 -5.275 ;
        RECT 16.155 -5.605 16.485 -5.275 ;
        RECT 14.795 -5.605 15.125 -5.275 ;
        RECT 13.435 -5.605 13.765 -5.275 ;
        RECT 12.075 -5.605 12.405 -5.275 ;
        RECT 10.715 -5.605 11.045 -5.275 ;
        RECT 9.355 -5.605 9.685 -5.275 ;
        RECT 7.995 -5.605 8.325 -5.275 ;
        RECT 6.635 -5.605 6.965 -5.275 ;
        RECT 5.275 -5.605 5.605 -5.275 ;
        RECT 3.915 -5.605 4.245 -5.275 ;
        RECT 2.555 -5.605 2.885 -5.275 ;
        RECT 1.195 -5.605 1.525 -5.275 ;
        RECT -0.165 -5.605 0.165 -5.275 ;
        RECT -1.525 -5.605 -1.195 -5.275 ;
        RECT -1.525 -5.6 678.475 -5.28 ;
        RECT 677.115 -5.605 677.445 -5.275 ;
        RECT 675.755 -5.605 676.085 -5.275 ;
        RECT 674.395 -5.605 674.725 -5.275 ;
        RECT 673.035 -5.605 673.365 -5.275 ;
        RECT 671.675 -5.605 672.005 -5.275 ;
        RECT 670.315 -5.605 670.645 -5.275 ;
        RECT 668.955 -5.605 669.285 -5.275 ;
        RECT 667.595 -5.605 667.925 -5.275 ;
        RECT 666.235 -5.605 666.565 -5.275 ;
        RECT 664.875 -5.605 665.205 -5.275 ;
        RECT 663.515 -5.605 663.845 -5.275 ;
        RECT 662.155 -5.605 662.485 -5.275 ;
        RECT 660.795 -5.605 661.125 -5.275 ;
        RECT 659.435 -5.605 659.765 -5.275 ;
        RECT 658.075 -5.605 658.405 -5.275 ;
        RECT 656.715 -5.605 657.045 -5.275 ;
        RECT 655.355 -5.605 655.685 -5.275 ;
        RECT 954.555 -5.605 954.885 -5.275 ;
        RECT 678.475 -5.6 954.885 -5.28 ;
        RECT 953.195 -5.605 953.525 -5.275 ;
        RECT 951.835 -5.605 952.165 -5.275 ;
        RECT 950.475 -5.605 950.805 -5.275 ;
        RECT 949.115 -5.605 949.445 -5.275 ;
        RECT 947.755 -5.605 948.085 -5.275 ;
        RECT 946.395 -5.605 946.725 -5.275 ;
        RECT 945.035 -5.605 945.365 -5.275 ;
        RECT 943.675 -5.605 944.005 -5.275 ;
        RECT 942.315 -5.605 942.645 -5.275 ;
        RECT 940.955 -5.605 941.285 -5.275 ;
        RECT 939.595 -5.605 939.925 -5.275 ;
        RECT 938.235 -5.605 938.565 -5.275 ;
        RECT 936.875 -5.605 937.205 -5.275 ;
        RECT 935.515 -5.605 935.845 -5.275 ;
        RECT 934.155 -5.605 934.485 -5.275 ;
        RECT 932.795 -5.605 933.125 -5.275 ;
        RECT 931.435 -5.605 931.765 -5.275 ;
        RECT 930.075 -5.605 930.405 -5.275 ;
        RECT 928.715 -5.605 929.045 -5.275 ;
        RECT 927.355 -5.605 927.685 -5.275 ;
        RECT 925.995 -5.605 926.325 -5.275 ;
        RECT 924.635 -5.605 924.965 -5.275 ;
        RECT 923.275 -5.605 923.605 -5.275 ;
        RECT 921.915 -5.605 922.245 -5.275 ;
        RECT 920.555 -5.605 920.885 -5.275 ;
        RECT 919.195 -5.605 919.525 -5.275 ;
        RECT 917.835 -5.605 918.165 -5.275 ;
        RECT 916.475 -5.605 916.805 -5.275 ;
        RECT 915.115 -5.605 915.445 -5.275 ;
        RECT 913.755 -5.605 914.085 -5.275 ;
        RECT 912.395 -5.605 912.725 -5.275 ;
        RECT 911.035 -5.605 911.365 -5.275 ;
        RECT 909.675 -5.605 910.005 -5.275 ;
        RECT 908.315 -5.605 908.645 -5.275 ;
        RECT 906.955 -5.605 907.285 -5.275 ;
        RECT 905.595 -5.605 905.925 -5.275 ;
        RECT 904.235 -5.605 904.565 -5.275 ;
        RECT 902.875 -5.605 903.205 -5.275 ;
        RECT 901.515 -5.605 901.845 -5.275 ;
        RECT 900.155 -5.605 900.485 -5.275 ;
        RECT 898.795 -5.605 899.125 -5.275 ;
        RECT 897.435 -5.605 897.765 -5.275 ;
        RECT 896.075 -5.605 896.405 -5.275 ;
        RECT 894.715 -5.605 895.045 -5.275 ;
        RECT 893.355 -5.605 893.685 -5.275 ;
        RECT 891.995 -5.605 892.325 -5.275 ;
        RECT 890.635 -5.605 890.965 -5.275 ;
        RECT 889.275 -5.605 889.605 -5.275 ;
        RECT 887.915 -5.605 888.245 -5.275 ;
        RECT 886.555 -5.605 886.885 -5.275 ;
        RECT 885.195 -5.605 885.525 -5.275 ;
        RECT 883.835 -5.605 884.165 -5.275 ;
        RECT 882.475 -5.605 882.805 -5.275 ;
        RECT 881.115 -5.605 881.445 -5.275 ;
        RECT 879.755 -5.605 880.085 -5.275 ;
        RECT 878.395 -5.605 878.725 -5.275 ;
        RECT 877.035 -5.605 877.365 -5.275 ;
        RECT 875.675 -5.605 876.005 -5.275 ;
        RECT 874.315 -5.605 874.645 -5.275 ;
        RECT 872.955 -5.605 873.285 -5.275 ;
        RECT 871.595 -5.605 871.925 -5.275 ;
        RECT 870.235 -5.605 870.565 -5.275 ;
        RECT 868.875 -5.605 869.205 -5.275 ;
        RECT 867.515 -5.605 867.845 -5.275 ;
        RECT 866.155 -5.605 866.485 -5.275 ;
        RECT 864.795 -5.605 865.125 -5.275 ;
        RECT 863.435 -5.605 863.765 -5.275 ;
        RECT 862.075 -5.605 862.405 -5.275 ;
        RECT 860.715 -5.605 861.045 -5.275 ;
        RECT 859.355 -5.605 859.685 -5.275 ;
        RECT 857.995 -5.605 858.325 -5.275 ;
        RECT 856.635 -5.605 856.965 -5.275 ;
        RECT 855.275 -5.605 855.605 -5.275 ;
        RECT 853.915 -5.605 854.245 -5.275 ;
        RECT 852.555 -5.605 852.885 -5.275 ;
        RECT 851.195 -5.605 851.525 -5.275 ;
        RECT 849.835 -5.605 850.165 -5.275 ;
        RECT 848.475 -5.605 848.805 -5.275 ;
        RECT 847.115 -5.605 847.445 -5.275 ;
        RECT 845.755 -5.605 846.085 -5.275 ;
        RECT 844.395 -5.605 844.725 -5.275 ;
        RECT 843.035 -5.605 843.365 -5.275 ;
        RECT 841.675 -5.605 842.005 -5.275 ;
        RECT 840.315 -5.605 840.645 -5.275 ;
        RECT 838.955 -5.605 839.285 -5.275 ;
        RECT 837.595 -5.605 837.925 -5.275 ;
        RECT 836.235 -5.605 836.565 -5.275 ;
        RECT 834.875 -5.605 835.205 -5.275 ;
        RECT 833.515 -5.605 833.845 -5.275 ;
        RECT 832.155 -5.605 832.485 -5.275 ;
        RECT 830.795 -5.605 831.125 -5.275 ;
        RECT 829.435 -5.605 829.765 -5.275 ;
        RECT 828.075 -5.605 828.405 -5.275 ;
        RECT 826.715 -5.605 827.045 -5.275 ;
        RECT 825.355 -5.605 825.685 -5.275 ;
        RECT 823.995 -5.605 824.325 -5.275 ;
        RECT 822.635 -5.605 822.965 -5.275 ;
        RECT 821.275 -5.605 821.605 -5.275 ;
        RECT 819.915 -5.605 820.245 -5.275 ;
        RECT 818.555 -5.605 818.885 -5.275 ;
        RECT 817.195 -5.605 817.525 -5.275 ;
        RECT 815.835 -5.605 816.165 -5.275 ;
        RECT 814.475 -5.605 814.805 -5.275 ;
        RECT 813.115 -5.605 813.445 -5.275 ;
        RECT 811.755 -5.605 812.085 -5.275 ;
        RECT 810.395 -5.605 810.725 -5.275 ;
        RECT 809.035 -5.605 809.365 -5.275 ;
        RECT 807.675 -5.605 808.005 -5.275 ;
        RECT 806.315 -5.605 806.645 -5.275 ;
        RECT 804.955 -5.605 805.285 -5.275 ;
        RECT 803.595 -5.605 803.925 -5.275 ;
        RECT 802.235 -5.605 802.565 -5.275 ;
        RECT 800.875 -5.605 801.205 -5.275 ;
        RECT 799.515 -5.605 799.845 -5.275 ;
        RECT 798.155 -5.605 798.485 -5.275 ;
        RECT 796.795 -5.605 797.125 -5.275 ;
        RECT 795.435 -5.605 795.765 -5.275 ;
        RECT 794.075 -5.605 794.405 -5.275 ;
        RECT 792.715 -5.605 793.045 -5.275 ;
        RECT 791.355 -5.605 791.685 -5.275 ;
        RECT 789.995 -5.605 790.325 -5.275 ;
        RECT 788.635 -5.605 788.965 -5.275 ;
        RECT 787.275 -5.605 787.605 -5.275 ;
        RECT 785.915 -5.605 786.245 -5.275 ;
        RECT 784.555 -5.605 784.885 -5.275 ;
        RECT 783.195 -5.605 783.525 -5.275 ;
        RECT 781.835 -5.605 782.165 -5.275 ;
        RECT 780.475 -5.605 780.805 -5.275 ;
        RECT 779.115 -5.605 779.445 -5.275 ;
        RECT 777.755 -5.605 778.085 -5.275 ;
        RECT 776.395 -5.605 776.725 -5.275 ;
        RECT 775.035 -5.605 775.365 -5.275 ;
        RECT 773.675 -5.605 774.005 -5.275 ;
        RECT 772.315 -5.605 772.645 -5.275 ;
        RECT 770.955 -5.605 771.285 -5.275 ;
        RECT 769.595 -5.605 769.925 -5.275 ;
        RECT 768.235 -5.605 768.565 -5.275 ;
        RECT 766.875 -5.605 767.205 -5.275 ;
        RECT 765.515 -5.605 765.845 -5.275 ;
        RECT 764.155 -5.605 764.485 -5.275 ;
        RECT 762.795 -5.605 763.125 -5.275 ;
        RECT 761.435 -5.605 761.765 -5.275 ;
        RECT 760.075 -5.605 760.405 -5.275 ;
        RECT 758.715 -5.605 759.045 -5.275 ;
        RECT 757.355 -5.605 757.685 -5.275 ;
        RECT 755.995 -5.605 756.325 -5.275 ;
        RECT 754.635 -5.605 754.965 -5.275 ;
        RECT 753.275 -5.605 753.605 -5.275 ;
        RECT 751.915 -5.605 752.245 -5.275 ;
        RECT 750.555 -5.605 750.885 -5.275 ;
        RECT 749.195 -5.605 749.525 -5.275 ;
        RECT 747.835 -5.605 748.165 -5.275 ;
        RECT 746.475 -5.605 746.805 -5.275 ;
        RECT 745.115 -5.605 745.445 -5.275 ;
        RECT 743.755 -5.605 744.085 -5.275 ;
        RECT 742.395 -5.605 742.725 -5.275 ;
        RECT 741.035 -5.605 741.365 -5.275 ;
        RECT 739.675 -5.605 740.005 -5.275 ;
        RECT 738.315 -5.605 738.645 -5.275 ;
        RECT 736.955 -5.605 737.285 -5.275 ;
        RECT 735.595 -5.605 735.925 -5.275 ;
        RECT 734.235 -5.605 734.565 -5.275 ;
        RECT 732.875 -5.605 733.205 -5.275 ;
        RECT 731.515 -5.605 731.845 -5.275 ;
        RECT 730.155 -5.605 730.485 -5.275 ;
        RECT 728.795 -5.605 729.125 -5.275 ;
        RECT 727.435 -5.605 727.765 -5.275 ;
        RECT 726.075 -5.605 726.405 -5.275 ;
        RECT 724.715 -5.605 725.045 -5.275 ;
        RECT 723.355 -5.605 723.685 -5.275 ;
        RECT 721.995 -5.605 722.325 -5.275 ;
        RECT 720.635 -5.605 720.965 -5.275 ;
        RECT 719.275 -5.605 719.605 -5.275 ;
        RECT 717.915 -5.605 718.245 -5.275 ;
        RECT 716.555 -5.605 716.885 -5.275 ;
        RECT 715.195 -5.605 715.525 -5.275 ;
        RECT 713.835 -5.605 714.165 -5.275 ;
        RECT 712.475 -5.605 712.805 -5.275 ;
        RECT 711.115 -5.605 711.445 -5.275 ;
        RECT 709.755 -5.605 710.085 -5.275 ;
        RECT 708.395 -5.605 708.725 -5.275 ;
        RECT 707.035 -5.605 707.365 -5.275 ;
        RECT 705.675 -5.605 706.005 -5.275 ;
        RECT 704.315 -5.605 704.645 -5.275 ;
        RECT 702.955 -5.605 703.285 -5.275 ;
        RECT 701.595 -5.605 701.925 -5.275 ;
        RECT 700.235 -5.605 700.565 -5.275 ;
        RECT 698.875 -5.605 699.205 -5.275 ;
        RECT 697.515 -5.605 697.845 -5.275 ;
        RECT 696.155 -5.605 696.485 -5.275 ;
        RECT 694.795 -5.605 695.125 -5.275 ;
        RECT 693.435 -5.605 693.765 -5.275 ;
        RECT 692.075 -5.605 692.405 -5.275 ;
        RECT 690.715 -5.605 691.045 -5.275 ;
        RECT 689.355 -5.605 689.685 -5.275 ;
        RECT 687.995 -5.605 688.325 -5.275 ;
        RECT 686.635 -5.605 686.965 -5.275 ;
        RECT 685.275 -5.605 685.605 -5.275 ;
        RECT 683.915 -5.605 684.245 -5.275 ;
        RECT 682.555 -5.605 682.885 -5.275 ;
        RECT 681.195 -5.605 681.525 -5.275 ;
        RECT 679.835 -5.605 680.165 -5.275 ;
        RECT 678.475 -5.605 678.805 -5.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -1.52 678.475 -1.2 ;
        RECT 677.115 -1.525 677.445 -1.195 ;
        RECT 675.755 -1.525 676.085 -1.195 ;
        RECT 674.395 -1.525 674.725 -1.195 ;
        RECT 673.035 -1.525 673.365 -1.195 ;
        RECT 671.675 -1.525 672.005 -1.195 ;
        RECT 670.315 -1.525 670.645 -1.195 ;
        RECT 668.955 -1.525 669.285 -1.195 ;
        RECT 667.595 -1.525 667.925 -1.195 ;
        RECT 666.235 -1.525 666.565 -1.195 ;
        RECT 664.875 -1.525 665.205 -1.195 ;
        RECT 663.515 -1.525 663.845 -1.195 ;
        RECT 662.155 -1.525 662.485 -1.195 ;
        RECT 660.795 -1.525 661.125 -1.195 ;
        RECT 659.435 -1.525 659.765 -1.195 ;
        RECT 658.075 -1.525 658.405 -1.195 ;
        RECT 656.715 -1.525 657.045 -1.195 ;
        RECT 655.355 -1.525 655.685 -1.195 ;
        RECT 653.995 -1.525 654.325 -1.195 ;
        RECT 652.635 -1.525 652.965 -1.195 ;
        RECT 651.275 -1.525 651.605 -1.195 ;
        RECT 649.915 -1.525 650.245 -1.195 ;
        RECT 648.555 -1.525 648.885 -1.195 ;
        RECT 647.195 -1.525 647.525 -1.195 ;
        RECT 645.835 -1.525 646.165 -1.195 ;
        RECT 644.475 -1.525 644.805 -1.195 ;
        RECT 643.115 -1.525 643.445 -1.195 ;
        RECT 641.755 -1.525 642.085 -1.195 ;
        RECT 640.395 -1.525 640.725 -1.195 ;
        RECT 639.035 -1.525 639.365 -1.195 ;
        RECT 637.675 -1.525 638.005 -1.195 ;
        RECT 636.315 -1.525 636.645 -1.195 ;
        RECT 634.955 -1.525 635.285 -1.195 ;
        RECT 633.595 -1.525 633.925 -1.195 ;
        RECT 632.235 -1.525 632.565 -1.195 ;
        RECT 630.875 -1.525 631.205 -1.195 ;
        RECT 629.515 -1.525 629.845 -1.195 ;
        RECT 628.155 -1.525 628.485 -1.195 ;
        RECT 626.795 -1.525 627.125 -1.195 ;
        RECT 625.435 -1.525 625.765 -1.195 ;
        RECT 624.075 -1.525 624.405 -1.195 ;
        RECT 622.715 -1.525 623.045 -1.195 ;
        RECT 621.355 -1.525 621.685 -1.195 ;
        RECT 619.995 -1.525 620.325 -1.195 ;
        RECT 618.635 -1.525 618.965 -1.195 ;
        RECT 617.275 -1.525 617.605 -1.195 ;
        RECT 615.915 -1.525 616.245 -1.195 ;
        RECT 614.555 -1.525 614.885 -1.195 ;
        RECT 613.195 -1.525 613.525 -1.195 ;
        RECT 611.835 -1.525 612.165 -1.195 ;
        RECT 610.475 -1.525 610.805 -1.195 ;
        RECT 609.115 -1.525 609.445 -1.195 ;
        RECT 607.755 -1.525 608.085 -1.195 ;
        RECT 606.395 -1.525 606.725 -1.195 ;
        RECT 605.035 -1.525 605.365 -1.195 ;
        RECT 603.675 -1.525 604.005 -1.195 ;
        RECT 602.315 -1.525 602.645 -1.195 ;
        RECT 600.955 -1.525 601.285 -1.195 ;
        RECT 599.595 -1.525 599.925 -1.195 ;
        RECT 598.235 -1.525 598.565 -1.195 ;
        RECT 596.875 -1.525 597.205 -1.195 ;
        RECT 595.515 -1.525 595.845 -1.195 ;
        RECT 594.155 -1.525 594.485 -1.195 ;
        RECT 592.795 -1.525 593.125 -1.195 ;
        RECT 591.435 -1.525 591.765 -1.195 ;
        RECT 590.075 -1.525 590.405 -1.195 ;
        RECT 588.715 -1.525 589.045 -1.195 ;
        RECT 587.355 -1.525 587.685 -1.195 ;
        RECT 585.995 -1.525 586.325 -1.195 ;
        RECT 584.635 -1.525 584.965 -1.195 ;
        RECT 583.275 -1.525 583.605 -1.195 ;
        RECT 581.915 -1.525 582.245 -1.195 ;
        RECT 580.555 -1.525 580.885 -1.195 ;
        RECT 579.195 -1.525 579.525 -1.195 ;
        RECT 577.835 -1.525 578.165 -1.195 ;
        RECT 576.475 -1.525 576.805 -1.195 ;
        RECT 575.115 -1.525 575.445 -1.195 ;
        RECT 573.755 -1.525 574.085 -1.195 ;
        RECT 572.395 -1.525 572.725 -1.195 ;
        RECT 571.035 -1.525 571.365 -1.195 ;
        RECT 569.675 -1.525 570.005 -1.195 ;
        RECT 568.315 -1.525 568.645 -1.195 ;
        RECT 566.955 -1.525 567.285 -1.195 ;
        RECT 565.595 -1.525 565.925 -1.195 ;
        RECT 564.235 -1.525 564.565 -1.195 ;
        RECT 562.875 -1.525 563.205 -1.195 ;
        RECT 561.515 -1.525 561.845 -1.195 ;
        RECT 560.155 -1.525 560.485 -1.195 ;
        RECT 558.795 -1.525 559.125 -1.195 ;
        RECT 557.435 -1.525 557.765 -1.195 ;
        RECT 556.075 -1.525 556.405 -1.195 ;
        RECT 554.715 -1.525 555.045 -1.195 ;
        RECT 553.355 -1.525 553.685 -1.195 ;
        RECT 551.995 -1.525 552.325 -1.195 ;
        RECT 550.635 -1.525 550.965 -1.195 ;
        RECT 549.275 -1.525 549.605 -1.195 ;
        RECT 547.915 -1.525 548.245 -1.195 ;
        RECT 546.555 -1.525 546.885 -1.195 ;
        RECT 545.195 -1.525 545.525 -1.195 ;
        RECT 543.835 -1.525 544.165 -1.195 ;
        RECT 542.475 -1.525 542.805 -1.195 ;
        RECT 541.115 -1.525 541.445 -1.195 ;
        RECT 539.755 -1.525 540.085 -1.195 ;
        RECT 538.395 -1.525 538.725 -1.195 ;
        RECT 537.035 -1.525 537.365 -1.195 ;
        RECT 535.675 -1.525 536.005 -1.195 ;
        RECT 534.315 -1.525 534.645 -1.195 ;
        RECT 532.955 -1.525 533.285 -1.195 ;
        RECT 531.595 -1.525 531.925 -1.195 ;
        RECT 530.235 -1.525 530.565 -1.195 ;
        RECT 528.875 -1.525 529.205 -1.195 ;
        RECT 527.515 -1.525 527.845 -1.195 ;
        RECT 526.155 -1.525 526.485 -1.195 ;
        RECT 524.795 -1.525 525.125 -1.195 ;
        RECT 523.435 -1.525 523.765 -1.195 ;
        RECT 522.075 -1.525 522.405 -1.195 ;
        RECT 520.715 -1.525 521.045 -1.195 ;
        RECT 519.355 -1.525 519.685 -1.195 ;
        RECT 517.995 -1.525 518.325 -1.195 ;
        RECT 516.635 -1.525 516.965 -1.195 ;
        RECT 515.275 -1.525 515.605 -1.195 ;
        RECT 513.915 -1.525 514.245 -1.195 ;
        RECT 512.555 -1.525 512.885 -1.195 ;
        RECT 511.195 -1.525 511.525 -1.195 ;
        RECT 509.835 -1.525 510.165 -1.195 ;
        RECT 508.475 -1.525 508.805 -1.195 ;
        RECT 507.115 -1.525 507.445 -1.195 ;
        RECT 505.755 -1.525 506.085 -1.195 ;
        RECT 504.395 -1.525 504.725 -1.195 ;
        RECT 503.035 -1.525 503.365 -1.195 ;
        RECT 501.675 -1.525 502.005 -1.195 ;
        RECT 500.315 -1.525 500.645 -1.195 ;
        RECT 498.955 -1.525 499.285 -1.195 ;
        RECT 497.595 -1.525 497.925 -1.195 ;
        RECT 496.235 -1.525 496.565 -1.195 ;
        RECT 494.875 -1.525 495.205 -1.195 ;
        RECT 493.515 -1.525 493.845 -1.195 ;
        RECT 492.155 -1.525 492.485 -1.195 ;
        RECT 490.795 -1.525 491.125 -1.195 ;
        RECT 489.435 -1.525 489.765 -1.195 ;
        RECT 488.075 -1.525 488.405 -1.195 ;
        RECT 486.715 -1.525 487.045 -1.195 ;
        RECT 485.355 -1.525 485.685 -1.195 ;
        RECT 483.995 -1.525 484.325 -1.195 ;
        RECT 482.635 -1.525 482.965 -1.195 ;
        RECT 481.275 -1.525 481.605 -1.195 ;
        RECT 479.915 -1.525 480.245 -1.195 ;
        RECT 478.555 -1.525 478.885 -1.195 ;
        RECT 477.195 -1.525 477.525 -1.195 ;
        RECT 475.835 -1.525 476.165 -1.195 ;
        RECT 474.475 -1.525 474.805 -1.195 ;
        RECT 473.115 -1.525 473.445 -1.195 ;
        RECT 471.755 -1.525 472.085 -1.195 ;
        RECT 470.395 -1.525 470.725 -1.195 ;
        RECT 469.035 -1.525 469.365 -1.195 ;
        RECT 467.675 -1.525 468.005 -1.195 ;
        RECT 466.315 -1.525 466.645 -1.195 ;
        RECT 464.955 -1.525 465.285 -1.195 ;
        RECT 463.595 -1.525 463.925 -1.195 ;
        RECT 462.235 -1.525 462.565 -1.195 ;
        RECT 460.875 -1.525 461.205 -1.195 ;
        RECT 459.515 -1.525 459.845 -1.195 ;
        RECT 458.155 -1.525 458.485 -1.195 ;
        RECT 456.795 -1.525 457.125 -1.195 ;
        RECT 455.435 -1.525 455.765 -1.195 ;
        RECT 454.075 -1.525 454.405 -1.195 ;
        RECT 452.715 -1.525 453.045 -1.195 ;
        RECT 451.355 -1.525 451.685 -1.195 ;
        RECT 449.995 -1.525 450.325 -1.195 ;
        RECT 448.635 -1.525 448.965 -1.195 ;
        RECT 447.275 -1.525 447.605 -1.195 ;
        RECT 445.915 -1.525 446.245 -1.195 ;
        RECT 444.555 -1.525 444.885 -1.195 ;
        RECT 443.195 -1.525 443.525 -1.195 ;
        RECT 441.835 -1.525 442.165 -1.195 ;
        RECT 440.475 -1.525 440.805 -1.195 ;
        RECT 439.115 -1.525 439.445 -1.195 ;
        RECT 437.755 -1.525 438.085 -1.195 ;
        RECT 436.395 -1.525 436.725 -1.195 ;
        RECT 435.035 -1.525 435.365 -1.195 ;
        RECT 433.675 -1.525 434.005 -1.195 ;
        RECT 432.315 -1.525 432.645 -1.195 ;
        RECT 430.955 -1.525 431.285 -1.195 ;
        RECT 429.595 -1.525 429.925 -1.195 ;
        RECT 428.235 -1.525 428.565 -1.195 ;
        RECT 426.875 -1.525 427.205 -1.195 ;
        RECT 425.515 -1.525 425.845 -1.195 ;
        RECT 424.155 -1.525 424.485 -1.195 ;
        RECT 422.795 -1.525 423.125 -1.195 ;
        RECT 421.435 -1.525 421.765 -1.195 ;
        RECT 420.075 -1.525 420.405 -1.195 ;
        RECT 418.715 -1.525 419.045 -1.195 ;
        RECT 417.355 -1.525 417.685 -1.195 ;
        RECT 415.995 -1.525 416.325 -1.195 ;
        RECT 414.635 -1.525 414.965 -1.195 ;
        RECT 413.275 -1.525 413.605 -1.195 ;
        RECT 411.915 -1.525 412.245 -1.195 ;
        RECT 410.555 -1.525 410.885 -1.195 ;
        RECT 409.195 -1.525 409.525 -1.195 ;
        RECT 407.835 -1.525 408.165 -1.195 ;
        RECT 406.475 -1.525 406.805 -1.195 ;
        RECT 405.115 -1.525 405.445 -1.195 ;
        RECT 403.755 -1.525 404.085 -1.195 ;
        RECT 402.395 -1.525 402.725 -1.195 ;
        RECT 401.035 -1.525 401.365 -1.195 ;
        RECT 399.675 -1.525 400.005 -1.195 ;
        RECT 398.315 -1.525 398.645 -1.195 ;
        RECT 396.955 -1.525 397.285 -1.195 ;
        RECT 395.595 -1.525 395.925 -1.195 ;
        RECT 394.235 -1.525 394.565 -1.195 ;
        RECT 392.875 -1.525 393.205 -1.195 ;
        RECT 391.515 -1.525 391.845 -1.195 ;
        RECT 390.155 -1.525 390.485 -1.195 ;
        RECT 388.795 -1.525 389.125 -1.195 ;
        RECT 387.435 -1.525 387.765 -1.195 ;
        RECT 386.075 -1.525 386.405 -1.195 ;
        RECT 384.715 -1.525 385.045 -1.195 ;
        RECT 383.355 -1.525 383.685 -1.195 ;
        RECT 381.995 -1.525 382.325 -1.195 ;
        RECT 380.635 -1.525 380.965 -1.195 ;
        RECT 379.275 -1.525 379.605 -1.195 ;
        RECT 377.915 -1.525 378.245 -1.195 ;
        RECT 376.555 -1.525 376.885 -1.195 ;
        RECT 375.195 -1.525 375.525 -1.195 ;
        RECT 373.835 -1.525 374.165 -1.195 ;
        RECT 372.475 -1.525 372.805 -1.195 ;
        RECT 371.115 -1.525 371.445 -1.195 ;
        RECT 369.755 -1.525 370.085 -1.195 ;
        RECT 368.395 -1.525 368.725 -1.195 ;
        RECT 367.035 -1.525 367.365 -1.195 ;
        RECT 365.675 -1.525 366.005 -1.195 ;
        RECT 364.315 -1.525 364.645 -1.195 ;
        RECT 362.955 -1.525 363.285 -1.195 ;
        RECT 361.595 -1.525 361.925 -1.195 ;
        RECT 360.235 -1.525 360.565 -1.195 ;
        RECT 358.875 -1.525 359.205 -1.195 ;
        RECT 357.515 -1.525 357.845 -1.195 ;
        RECT 356.155 -1.525 356.485 -1.195 ;
        RECT 354.795 -1.525 355.125 -1.195 ;
        RECT 353.435 -1.525 353.765 -1.195 ;
        RECT 352.075 -1.525 352.405 -1.195 ;
        RECT 350.715 -1.525 351.045 -1.195 ;
        RECT 349.355 -1.525 349.685 -1.195 ;
        RECT 347.995 -1.525 348.325 -1.195 ;
        RECT 346.635 -1.525 346.965 -1.195 ;
        RECT 345.275 -1.525 345.605 -1.195 ;
        RECT 343.915 -1.525 344.245 -1.195 ;
        RECT 342.555 -1.525 342.885 -1.195 ;
        RECT 341.195 -1.525 341.525 -1.195 ;
        RECT 339.835 -1.525 340.165 -1.195 ;
        RECT 338.475 -1.525 338.805 -1.195 ;
        RECT 337.115 -1.525 337.445 -1.195 ;
        RECT 335.755 -1.525 336.085 -1.195 ;
        RECT 334.395 -1.525 334.725 -1.195 ;
        RECT 333.035 -1.525 333.365 -1.195 ;
        RECT 331.675 -1.525 332.005 -1.195 ;
        RECT 330.315 -1.525 330.645 -1.195 ;
        RECT 328.955 -1.525 329.285 -1.195 ;
        RECT 327.595 -1.525 327.925 -1.195 ;
        RECT 326.235 -1.525 326.565 -1.195 ;
        RECT 324.875 -1.525 325.205 -1.195 ;
        RECT 323.515 -1.525 323.845 -1.195 ;
        RECT 322.155 -1.525 322.485 -1.195 ;
        RECT 320.795 -1.525 321.125 -1.195 ;
        RECT 319.435 -1.525 319.765 -1.195 ;
        RECT 318.075 -1.525 318.405 -1.195 ;
        RECT 316.715 -1.525 317.045 -1.195 ;
        RECT 315.355 -1.525 315.685 -1.195 ;
        RECT 313.995 -1.525 314.325 -1.195 ;
        RECT 312.635 -1.525 312.965 -1.195 ;
        RECT 311.275 -1.525 311.605 -1.195 ;
        RECT 309.915 -1.525 310.245 -1.195 ;
        RECT 308.555 -1.525 308.885 -1.195 ;
        RECT 307.195 -1.525 307.525 -1.195 ;
        RECT 305.835 -1.525 306.165 -1.195 ;
        RECT 304.475 -1.525 304.805 -1.195 ;
        RECT 303.115 -1.525 303.445 -1.195 ;
        RECT 301.755 -1.525 302.085 -1.195 ;
        RECT 300.395 -1.525 300.725 -1.195 ;
        RECT 299.035 -1.525 299.365 -1.195 ;
        RECT 297.675 -1.525 298.005 -1.195 ;
        RECT 296.315 -1.525 296.645 -1.195 ;
        RECT 294.955 -1.525 295.285 -1.195 ;
        RECT 293.595 -1.525 293.925 -1.195 ;
        RECT 292.235 -1.525 292.565 -1.195 ;
        RECT 290.875 -1.525 291.205 -1.195 ;
        RECT 289.515 -1.525 289.845 -1.195 ;
        RECT 288.155 -1.525 288.485 -1.195 ;
        RECT 286.795 -1.525 287.125 -1.195 ;
        RECT 285.435 -1.525 285.765 -1.195 ;
        RECT 284.075 -1.525 284.405 -1.195 ;
        RECT 282.715 -1.525 283.045 -1.195 ;
        RECT 281.355 -1.525 281.685 -1.195 ;
        RECT 279.995 -1.525 280.325 -1.195 ;
        RECT 278.635 -1.525 278.965 -1.195 ;
        RECT 277.275 -1.525 277.605 -1.195 ;
        RECT 275.915 -1.525 276.245 -1.195 ;
        RECT 274.555 -1.525 274.885 -1.195 ;
        RECT 273.195 -1.525 273.525 -1.195 ;
        RECT 271.835 -1.525 272.165 -1.195 ;
        RECT 270.475 -1.525 270.805 -1.195 ;
        RECT 269.115 -1.525 269.445 -1.195 ;
        RECT 267.755 -1.525 268.085 -1.195 ;
        RECT 266.395 -1.525 266.725 -1.195 ;
        RECT 265.035 -1.525 265.365 -1.195 ;
        RECT 263.675 -1.525 264.005 -1.195 ;
        RECT 262.315 -1.525 262.645 -1.195 ;
        RECT 260.955 -1.525 261.285 -1.195 ;
        RECT 259.595 -1.525 259.925 -1.195 ;
        RECT 258.235 -1.525 258.565 -1.195 ;
        RECT 256.875 -1.525 257.205 -1.195 ;
        RECT 255.515 -1.525 255.845 -1.195 ;
        RECT 254.155 -1.525 254.485 -1.195 ;
        RECT 252.795 -1.525 253.125 -1.195 ;
        RECT 251.435 -1.525 251.765 -1.195 ;
        RECT 250.075 -1.525 250.405 -1.195 ;
        RECT 248.715 -1.525 249.045 -1.195 ;
        RECT 247.355 -1.525 247.685 -1.195 ;
        RECT 245.995 -1.525 246.325 -1.195 ;
        RECT 244.635 -1.525 244.965 -1.195 ;
        RECT 243.275 -1.525 243.605 -1.195 ;
        RECT 241.915 -1.525 242.245 -1.195 ;
        RECT 240.555 -1.525 240.885 -1.195 ;
        RECT 239.195 -1.525 239.525 -1.195 ;
        RECT 237.835 -1.525 238.165 -1.195 ;
        RECT 236.475 -1.525 236.805 -1.195 ;
        RECT 235.115 -1.525 235.445 -1.195 ;
        RECT 233.755 -1.525 234.085 -1.195 ;
        RECT 232.395 -1.525 232.725 -1.195 ;
        RECT 231.035 -1.525 231.365 -1.195 ;
        RECT 229.675 -1.525 230.005 -1.195 ;
        RECT 228.315 -1.525 228.645 -1.195 ;
        RECT 226.955 -1.525 227.285 -1.195 ;
        RECT 225.595 -1.525 225.925 -1.195 ;
        RECT 224.235 -1.525 224.565 -1.195 ;
        RECT 222.875 -1.525 223.205 -1.195 ;
        RECT 221.515 -1.525 221.845 -1.195 ;
        RECT 220.155 -1.525 220.485 -1.195 ;
        RECT 218.795 -1.525 219.125 -1.195 ;
        RECT 217.435 -1.525 217.765 -1.195 ;
        RECT 216.075 -1.525 216.405 -1.195 ;
        RECT 214.715 -1.525 215.045 -1.195 ;
        RECT 213.355 -1.525 213.685 -1.195 ;
        RECT 211.995 -1.525 212.325 -1.195 ;
        RECT 210.635 -1.525 210.965 -1.195 ;
        RECT 209.275 -1.525 209.605 -1.195 ;
        RECT 207.915 -1.525 208.245 -1.195 ;
        RECT 206.555 -1.525 206.885 -1.195 ;
        RECT 205.195 -1.525 205.525 -1.195 ;
        RECT 203.835 -1.525 204.165 -1.195 ;
        RECT 202.475 -1.525 202.805 -1.195 ;
        RECT 201.115 -1.525 201.445 -1.195 ;
        RECT 199.755 -1.525 200.085 -1.195 ;
        RECT 198.395 -1.525 198.725 -1.195 ;
        RECT 197.035 -1.525 197.365 -1.195 ;
        RECT 195.675 -1.525 196.005 -1.195 ;
        RECT 194.315 -1.525 194.645 -1.195 ;
        RECT 192.955 -1.525 193.285 -1.195 ;
        RECT 191.595 -1.525 191.925 -1.195 ;
        RECT 190.235 -1.525 190.565 -1.195 ;
        RECT 188.875 -1.525 189.205 -1.195 ;
        RECT 187.515 -1.525 187.845 -1.195 ;
        RECT 186.155 -1.525 186.485 -1.195 ;
        RECT 184.795 -1.525 185.125 -1.195 ;
        RECT 183.435 -1.525 183.765 -1.195 ;
        RECT 182.075 -1.525 182.405 -1.195 ;
        RECT 180.715 -1.525 181.045 -1.195 ;
        RECT 179.355 -1.525 179.685 -1.195 ;
        RECT 177.995 -1.525 178.325 -1.195 ;
        RECT 176.635 -1.525 176.965 -1.195 ;
        RECT 175.275 -1.525 175.605 -1.195 ;
        RECT 173.915 -1.525 174.245 -1.195 ;
        RECT 172.555 -1.525 172.885 -1.195 ;
        RECT 171.195 -1.525 171.525 -1.195 ;
        RECT 169.835 -1.525 170.165 -1.195 ;
        RECT 168.475 -1.525 168.805 -1.195 ;
        RECT 167.115 -1.525 167.445 -1.195 ;
        RECT 165.755 -1.525 166.085 -1.195 ;
        RECT 164.395 -1.525 164.725 -1.195 ;
        RECT 163.035 -1.525 163.365 -1.195 ;
        RECT 161.675 -1.525 162.005 -1.195 ;
        RECT 160.315 -1.525 160.645 -1.195 ;
        RECT 158.955 -1.525 159.285 -1.195 ;
        RECT 157.595 -1.525 157.925 -1.195 ;
        RECT 156.235 -1.525 156.565 -1.195 ;
        RECT 154.875 -1.525 155.205 -1.195 ;
        RECT 153.515 -1.525 153.845 -1.195 ;
        RECT 152.155 -1.525 152.485 -1.195 ;
        RECT 150.795 -1.525 151.125 -1.195 ;
        RECT 149.435 -1.525 149.765 -1.195 ;
        RECT 148.075 -1.525 148.405 -1.195 ;
        RECT 146.715 -1.525 147.045 -1.195 ;
        RECT 145.355 -1.525 145.685 -1.195 ;
        RECT 143.995 -1.525 144.325 -1.195 ;
        RECT 142.635 -1.525 142.965 -1.195 ;
        RECT 141.275 -1.525 141.605 -1.195 ;
        RECT 139.915 -1.525 140.245 -1.195 ;
        RECT 138.555 -1.525 138.885 -1.195 ;
        RECT 137.195 -1.525 137.525 -1.195 ;
        RECT 135.835 -1.525 136.165 -1.195 ;
        RECT 134.475 -1.525 134.805 -1.195 ;
        RECT 133.115 -1.525 133.445 -1.195 ;
        RECT 131.755 -1.525 132.085 -1.195 ;
        RECT 130.395 -1.525 130.725 -1.195 ;
        RECT 129.035 -1.525 129.365 -1.195 ;
        RECT 127.675 -1.525 128.005 -1.195 ;
        RECT 126.315 -1.525 126.645 -1.195 ;
        RECT 124.955 -1.525 125.285 -1.195 ;
        RECT 123.595 -1.525 123.925 -1.195 ;
        RECT 122.235 -1.525 122.565 -1.195 ;
        RECT 120.875 -1.525 121.205 -1.195 ;
        RECT 119.515 -1.525 119.845 -1.195 ;
        RECT 118.155 -1.525 118.485 -1.195 ;
        RECT 116.795 -1.525 117.125 -1.195 ;
        RECT 115.435 -1.525 115.765 -1.195 ;
        RECT 114.075 -1.525 114.405 -1.195 ;
        RECT 112.715 -1.525 113.045 -1.195 ;
        RECT 111.355 -1.525 111.685 -1.195 ;
        RECT 109.995 -1.525 110.325 -1.195 ;
        RECT 108.635 -1.525 108.965 -1.195 ;
        RECT 107.275 -1.525 107.605 -1.195 ;
        RECT 105.915 -1.525 106.245 -1.195 ;
        RECT 104.555 -1.525 104.885 -1.195 ;
        RECT 103.195 -1.525 103.525 -1.195 ;
        RECT 101.835 -1.525 102.165 -1.195 ;
        RECT 100.475 -1.525 100.805 -1.195 ;
        RECT 99.115 -1.525 99.445 -1.195 ;
        RECT 97.755 -1.525 98.085 -1.195 ;
        RECT 96.395 -1.525 96.725 -1.195 ;
        RECT 95.035 -1.525 95.365 -1.195 ;
        RECT 93.675 -1.525 94.005 -1.195 ;
        RECT 92.315 -1.525 92.645 -1.195 ;
        RECT 90.955 -1.525 91.285 -1.195 ;
        RECT 89.595 -1.525 89.925 -1.195 ;
        RECT 88.235 -1.525 88.565 -1.195 ;
        RECT 86.875 -1.525 87.205 -1.195 ;
        RECT 85.515 -1.525 85.845 -1.195 ;
        RECT 84.155 -1.525 84.485 -1.195 ;
        RECT 82.795 -1.525 83.125 -1.195 ;
        RECT 81.435 -1.525 81.765 -1.195 ;
        RECT 80.075 -1.525 80.405 -1.195 ;
        RECT 78.715 -1.525 79.045 -1.195 ;
        RECT 77.355 -1.525 77.685 -1.195 ;
        RECT 75.995 -1.525 76.325 -1.195 ;
        RECT 74.635 -1.525 74.965 -1.195 ;
        RECT 73.275 -1.525 73.605 -1.195 ;
        RECT 71.915 -1.525 72.245 -1.195 ;
        RECT 70.555 -1.525 70.885 -1.195 ;
        RECT 69.195 -1.525 69.525 -1.195 ;
        RECT 67.835 -1.525 68.165 -1.195 ;
        RECT 66.475 -1.525 66.805 -1.195 ;
        RECT 65.115 -1.525 65.445 -1.195 ;
        RECT 63.755 -1.525 64.085 -1.195 ;
        RECT 62.395 -1.525 62.725 -1.195 ;
        RECT 61.035 -1.525 61.365 -1.195 ;
        RECT 59.675 -1.525 60.005 -1.195 ;
        RECT 58.315 -1.525 58.645 -1.195 ;
        RECT 56.955 -1.525 57.285 -1.195 ;
        RECT 55.595 -1.525 55.925 -1.195 ;
        RECT 54.235 -1.525 54.565 -1.195 ;
        RECT 52.875 -1.525 53.205 -1.195 ;
        RECT 51.515 -1.525 51.845 -1.195 ;
        RECT 50.155 -1.525 50.485 -1.195 ;
        RECT 48.795 -1.525 49.125 -1.195 ;
        RECT 47.435 -1.525 47.765 -1.195 ;
        RECT 46.075 -1.525 46.405 -1.195 ;
        RECT 44.715 -1.525 45.045 -1.195 ;
        RECT 43.355 -1.525 43.685 -1.195 ;
        RECT 41.995 -1.525 42.325 -1.195 ;
        RECT 40.635 -1.525 40.965 -1.195 ;
        RECT 39.275 -1.525 39.605 -1.195 ;
        RECT 37.915 -1.525 38.245 -1.195 ;
        RECT 36.555 -1.525 36.885 -1.195 ;
        RECT 35.195 -1.525 35.525 -1.195 ;
        RECT 33.835 -1.525 34.165 -1.195 ;
        RECT 32.475 -1.525 32.805 -1.195 ;
        RECT 31.115 -1.525 31.445 -1.195 ;
        RECT 29.755 -1.525 30.085 -1.195 ;
        RECT 28.395 -1.525 28.725 -1.195 ;
        RECT 27.035 -1.525 27.365 -1.195 ;
        RECT 25.675 -1.525 26.005 -1.195 ;
        RECT 24.315 -1.525 24.645 -1.195 ;
        RECT 22.955 -1.525 23.285 -1.195 ;
        RECT 21.595 -1.525 21.925 -1.195 ;
        RECT 20.235 -1.525 20.565 -1.195 ;
        RECT 18.875 -1.525 19.205 -1.195 ;
        RECT 17.515 -1.525 17.845 -1.195 ;
        RECT 16.155 -1.525 16.485 -1.195 ;
        RECT 14.795 -1.525 15.125 -1.195 ;
        RECT 13.435 -1.525 13.765 -1.195 ;
        RECT 12.075 -1.525 12.405 -1.195 ;
        RECT 10.715 -1.525 11.045 -1.195 ;
        RECT 9.355 -1.525 9.685 -1.195 ;
        RECT 7.995 -1.525 8.325 -1.195 ;
        RECT 6.635 -1.525 6.965 -1.195 ;
        RECT 5.275 -1.525 5.605 -1.195 ;
        RECT 3.915 -1.525 4.245 -1.195 ;
        RECT 2.555 -1.525 2.885 -1.195 ;
        RECT 1.195 -1.525 1.525 -1.195 ;
        RECT -0.165 -1.525 0.165 -1.195 ;
        RECT -1.525 -1.525 -1.195 -1.195 ;
        RECT 954.555 -1.525 954.885 -1.195 ;
        RECT 678.475 -1.52 954.885 -1.2 ;
        RECT 953.195 -1.525 953.525 -1.195 ;
        RECT 951.835 -1.525 952.165 -1.195 ;
        RECT 950.475 -1.525 950.805 -1.195 ;
        RECT 949.115 -1.525 949.445 -1.195 ;
        RECT 947.755 -1.525 948.085 -1.195 ;
        RECT 946.395 -1.525 946.725 -1.195 ;
        RECT 945.035 -1.525 945.365 -1.195 ;
        RECT 943.675 -1.525 944.005 -1.195 ;
        RECT 942.315 -1.525 942.645 -1.195 ;
        RECT 940.955 -1.525 941.285 -1.195 ;
        RECT 939.595 -1.525 939.925 -1.195 ;
        RECT 938.235 -1.525 938.565 -1.195 ;
        RECT 936.875 -1.525 937.205 -1.195 ;
        RECT 935.515 -1.525 935.845 -1.195 ;
        RECT 934.155 -1.525 934.485 -1.195 ;
        RECT 932.795 -1.525 933.125 -1.195 ;
        RECT 931.435 -1.525 931.765 -1.195 ;
        RECT 930.075 -1.525 930.405 -1.195 ;
        RECT 928.715 -1.525 929.045 -1.195 ;
        RECT 927.355 -1.525 927.685 -1.195 ;
        RECT 925.995 -1.525 926.325 -1.195 ;
        RECT 924.635 -1.525 924.965 -1.195 ;
        RECT 923.275 -1.525 923.605 -1.195 ;
        RECT 921.915 -1.525 922.245 -1.195 ;
        RECT 920.555 -1.525 920.885 -1.195 ;
        RECT 919.195 -1.525 919.525 -1.195 ;
        RECT 917.835 -1.525 918.165 -1.195 ;
        RECT 916.475 -1.525 916.805 -1.195 ;
        RECT 915.115 -1.525 915.445 -1.195 ;
        RECT 913.755 -1.525 914.085 -1.195 ;
        RECT 912.395 -1.525 912.725 -1.195 ;
        RECT 911.035 -1.525 911.365 -1.195 ;
        RECT 909.675 -1.525 910.005 -1.195 ;
        RECT 908.315 -1.525 908.645 -1.195 ;
        RECT 906.955 -1.525 907.285 -1.195 ;
        RECT 905.595 -1.525 905.925 -1.195 ;
        RECT 904.235 -1.525 904.565 -1.195 ;
        RECT 902.875 -1.525 903.205 -1.195 ;
        RECT 901.515 -1.525 901.845 -1.195 ;
        RECT 900.155 -1.525 900.485 -1.195 ;
        RECT 898.795 -1.525 899.125 -1.195 ;
        RECT 897.435 -1.525 897.765 -1.195 ;
        RECT 896.075 -1.525 896.405 -1.195 ;
        RECT 894.715 -1.525 895.045 -1.195 ;
        RECT 893.355 -1.525 893.685 -1.195 ;
        RECT 891.995 -1.525 892.325 -1.195 ;
        RECT 890.635 -1.525 890.965 -1.195 ;
        RECT 889.275 -1.525 889.605 -1.195 ;
        RECT 887.915 -1.525 888.245 -1.195 ;
        RECT 886.555 -1.525 886.885 -1.195 ;
        RECT 885.195 -1.525 885.525 -1.195 ;
        RECT 883.835 -1.525 884.165 -1.195 ;
        RECT 882.475 -1.525 882.805 -1.195 ;
        RECT 881.115 -1.525 881.445 -1.195 ;
        RECT 879.755 -1.525 880.085 -1.195 ;
        RECT 878.395 -1.525 878.725 -1.195 ;
        RECT 877.035 -1.525 877.365 -1.195 ;
        RECT 875.675 -1.525 876.005 -1.195 ;
        RECT 874.315 -1.525 874.645 -1.195 ;
        RECT 872.955 -1.525 873.285 -1.195 ;
        RECT 871.595 -1.525 871.925 -1.195 ;
        RECT 870.235 -1.525 870.565 -1.195 ;
        RECT 868.875 -1.525 869.205 -1.195 ;
        RECT 867.515 -1.525 867.845 -1.195 ;
        RECT 866.155 -1.525 866.485 -1.195 ;
        RECT 864.795 -1.525 865.125 -1.195 ;
        RECT 863.435 -1.525 863.765 -1.195 ;
        RECT 862.075 -1.525 862.405 -1.195 ;
        RECT 860.715 -1.525 861.045 -1.195 ;
        RECT 859.355 -1.525 859.685 -1.195 ;
        RECT 857.995 -1.525 858.325 -1.195 ;
        RECT 856.635 -1.525 856.965 -1.195 ;
        RECT 855.275 -1.525 855.605 -1.195 ;
        RECT 853.915 -1.525 854.245 -1.195 ;
        RECT 852.555 -1.525 852.885 -1.195 ;
        RECT 851.195 -1.525 851.525 -1.195 ;
        RECT 849.835 -1.525 850.165 -1.195 ;
        RECT 848.475 -1.525 848.805 -1.195 ;
        RECT 847.115 -1.525 847.445 -1.195 ;
        RECT 845.755 -1.525 846.085 -1.195 ;
        RECT 844.395 -1.525 844.725 -1.195 ;
        RECT 843.035 -1.525 843.365 -1.195 ;
        RECT 841.675 -1.525 842.005 -1.195 ;
        RECT 840.315 -1.525 840.645 -1.195 ;
        RECT 838.955 -1.525 839.285 -1.195 ;
        RECT 837.595 -1.525 837.925 -1.195 ;
        RECT 836.235 -1.525 836.565 -1.195 ;
        RECT 834.875 -1.525 835.205 -1.195 ;
        RECT 833.515 -1.525 833.845 -1.195 ;
        RECT 832.155 -1.525 832.485 -1.195 ;
        RECT 830.795 -1.525 831.125 -1.195 ;
        RECT 829.435 -1.525 829.765 -1.195 ;
        RECT 828.075 -1.525 828.405 -1.195 ;
        RECT 826.715 -1.525 827.045 -1.195 ;
        RECT 825.355 -1.525 825.685 -1.195 ;
        RECT 823.995 -1.525 824.325 -1.195 ;
        RECT 822.635 -1.525 822.965 -1.195 ;
        RECT 821.275 -1.525 821.605 -1.195 ;
        RECT 819.915 -1.525 820.245 -1.195 ;
        RECT 818.555 -1.525 818.885 -1.195 ;
        RECT 817.195 -1.525 817.525 -1.195 ;
        RECT 815.835 -1.525 816.165 -1.195 ;
        RECT 814.475 -1.525 814.805 -1.195 ;
        RECT 813.115 -1.525 813.445 -1.195 ;
        RECT 811.755 -1.525 812.085 -1.195 ;
        RECT 810.395 -1.525 810.725 -1.195 ;
        RECT 809.035 -1.525 809.365 -1.195 ;
        RECT 807.675 -1.525 808.005 -1.195 ;
        RECT 806.315 -1.525 806.645 -1.195 ;
        RECT 804.955 -1.525 805.285 -1.195 ;
        RECT 803.595 -1.525 803.925 -1.195 ;
        RECT 802.235 -1.525 802.565 -1.195 ;
        RECT 800.875 -1.525 801.205 -1.195 ;
        RECT 799.515 -1.525 799.845 -1.195 ;
        RECT 798.155 -1.525 798.485 -1.195 ;
        RECT 796.795 -1.525 797.125 -1.195 ;
        RECT 795.435 -1.525 795.765 -1.195 ;
        RECT 794.075 -1.525 794.405 -1.195 ;
        RECT 792.715 -1.525 793.045 -1.195 ;
        RECT 791.355 -1.525 791.685 -1.195 ;
        RECT 789.995 -1.525 790.325 -1.195 ;
        RECT 788.635 -1.525 788.965 -1.195 ;
        RECT 787.275 -1.525 787.605 -1.195 ;
        RECT 785.915 -1.525 786.245 -1.195 ;
        RECT 784.555 -1.525 784.885 -1.195 ;
        RECT 783.195 -1.525 783.525 -1.195 ;
        RECT 781.835 -1.525 782.165 -1.195 ;
        RECT 780.475 -1.525 780.805 -1.195 ;
        RECT 779.115 -1.525 779.445 -1.195 ;
        RECT 777.755 -1.525 778.085 -1.195 ;
        RECT 776.395 -1.525 776.725 -1.195 ;
        RECT 775.035 -1.525 775.365 -1.195 ;
        RECT 773.675 -1.525 774.005 -1.195 ;
        RECT 772.315 -1.525 772.645 -1.195 ;
        RECT 770.955 -1.525 771.285 -1.195 ;
        RECT 769.595 -1.525 769.925 -1.195 ;
        RECT 768.235 -1.525 768.565 -1.195 ;
        RECT 766.875 -1.525 767.205 -1.195 ;
        RECT 765.515 -1.525 765.845 -1.195 ;
        RECT 764.155 -1.525 764.485 -1.195 ;
        RECT 762.795 -1.525 763.125 -1.195 ;
        RECT 761.435 -1.525 761.765 -1.195 ;
        RECT 760.075 -1.525 760.405 -1.195 ;
        RECT 758.715 -1.525 759.045 -1.195 ;
        RECT 757.355 -1.525 757.685 -1.195 ;
        RECT 755.995 -1.525 756.325 -1.195 ;
        RECT 754.635 -1.525 754.965 -1.195 ;
        RECT 753.275 -1.525 753.605 -1.195 ;
        RECT 751.915 -1.525 752.245 -1.195 ;
        RECT 750.555 -1.525 750.885 -1.195 ;
        RECT 749.195 -1.525 749.525 -1.195 ;
        RECT 747.835 -1.525 748.165 -1.195 ;
        RECT 746.475 -1.525 746.805 -1.195 ;
        RECT 745.115 -1.525 745.445 -1.195 ;
        RECT 743.755 -1.525 744.085 -1.195 ;
        RECT 742.395 -1.525 742.725 -1.195 ;
        RECT 741.035 -1.525 741.365 -1.195 ;
        RECT 739.675 -1.525 740.005 -1.195 ;
        RECT 738.315 -1.525 738.645 -1.195 ;
        RECT 736.955 -1.525 737.285 -1.195 ;
        RECT 735.595 -1.525 735.925 -1.195 ;
        RECT 734.235 -1.525 734.565 -1.195 ;
        RECT 732.875 -1.525 733.205 -1.195 ;
        RECT 731.515 -1.525 731.845 -1.195 ;
        RECT 730.155 -1.525 730.485 -1.195 ;
        RECT 728.795 -1.525 729.125 -1.195 ;
        RECT 727.435 -1.525 727.765 -1.195 ;
        RECT 726.075 -1.525 726.405 -1.195 ;
        RECT 724.715 -1.525 725.045 -1.195 ;
        RECT 723.355 -1.525 723.685 -1.195 ;
        RECT 721.995 -1.525 722.325 -1.195 ;
        RECT 720.635 -1.525 720.965 -1.195 ;
        RECT 719.275 -1.525 719.605 -1.195 ;
        RECT 717.915 -1.525 718.245 -1.195 ;
        RECT 716.555 -1.525 716.885 -1.195 ;
        RECT 715.195 -1.525 715.525 -1.195 ;
        RECT 713.835 -1.525 714.165 -1.195 ;
        RECT 712.475 -1.525 712.805 -1.195 ;
        RECT 711.115 -1.525 711.445 -1.195 ;
        RECT 709.755 -1.525 710.085 -1.195 ;
        RECT 708.395 -1.525 708.725 -1.195 ;
        RECT 707.035 -1.525 707.365 -1.195 ;
        RECT 705.675 -1.525 706.005 -1.195 ;
        RECT 704.315 -1.525 704.645 -1.195 ;
        RECT 702.955 -1.525 703.285 -1.195 ;
        RECT 701.595 -1.525 701.925 -1.195 ;
        RECT 700.235 -1.525 700.565 -1.195 ;
        RECT 698.875 -1.525 699.205 -1.195 ;
        RECT 697.515 -1.525 697.845 -1.195 ;
        RECT 696.155 -1.525 696.485 -1.195 ;
        RECT 694.795 -1.525 695.125 -1.195 ;
        RECT 693.435 -1.525 693.765 -1.195 ;
        RECT 692.075 -1.525 692.405 -1.195 ;
        RECT 690.715 -1.525 691.045 -1.195 ;
        RECT 689.355 -1.525 689.685 -1.195 ;
        RECT 687.995 -1.525 688.325 -1.195 ;
        RECT 686.635 -1.525 686.965 -1.195 ;
        RECT 685.275 -1.525 685.605 -1.195 ;
        RECT 683.915 -1.525 684.245 -1.195 ;
        RECT 682.555 -1.525 682.885 -1.195 ;
        RECT 681.195 -1.525 681.525 -1.195 ;
        RECT 679.835 -1.525 680.165 -1.195 ;
        RECT 678.475 -1.525 678.805 -1.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 656.715 -2.885 657.045 -2.555 ;
        RECT 655.355 -2.885 655.685 -2.555 ;
        RECT 653.995 -2.885 654.325 -2.555 ;
        RECT 652.635 -2.885 652.965 -2.555 ;
        RECT 651.275 -2.885 651.605 -2.555 ;
        RECT 649.915 -2.885 650.245 -2.555 ;
        RECT 648.555 -2.885 648.885 -2.555 ;
        RECT 647.195 -2.885 647.525 -2.555 ;
        RECT 645.835 -2.885 646.165 -2.555 ;
        RECT 644.475 -2.885 644.805 -2.555 ;
        RECT 643.115 -2.885 643.445 -2.555 ;
        RECT 641.755 -2.885 642.085 -2.555 ;
        RECT 640.395 -2.885 640.725 -2.555 ;
        RECT 639.035 -2.885 639.365 -2.555 ;
        RECT 637.675 -2.885 638.005 -2.555 ;
        RECT 636.315 -2.885 636.645 -2.555 ;
        RECT 634.955 -2.885 635.285 -2.555 ;
        RECT 633.595 -2.885 633.925 -2.555 ;
        RECT 632.235 -2.885 632.565 -2.555 ;
        RECT 630.875 -2.885 631.205 -2.555 ;
        RECT 629.515 -2.885 629.845 -2.555 ;
        RECT 628.155 -2.885 628.485 -2.555 ;
        RECT 626.795 -2.885 627.125 -2.555 ;
        RECT 625.435 -2.885 625.765 -2.555 ;
        RECT 624.075 -2.885 624.405 -2.555 ;
        RECT 622.715 -2.885 623.045 -2.555 ;
        RECT 621.355 -2.885 621.685 -2.555 ;
        RECT 619.995 -2.885 620.325 -2.555 ;
        RECT 618.635 -2.885 618.965 -2.555 ;
        RECT 617.275 -2.885 617.605 -2.555 ;
        RECT 615.915 -2.885 616.245 -2.555 ;
        RECT 614.555 -2.885 614.885 -2.555 ;
        RECT 613.195 -2.885 613.525 -2.555 ;
        RECT 611.835 -2.885 612.165 -2.555 ;
        RECT 610.475 -2.885 610.805 -2.555 ;
        RECT 609.115 -2.885 609.445 -2.555 ;
        RECT 607.755 -2.885 608.085 -2.555 ;
        RECT 606.395 -2.885 606.725 -2.555 ;
        RECT 605.035 -2.885 605.365 -2.555 ;
        RECT 603.675 -2.885 604.005 -2.555 ;
        RECT 602.315 -2.885 602.645 -2.555 ;
        RECT 600.955 -2.885 601.285 -2.555 ;
        RECT 599.595 -2.885 599.925 -2.555 ;
        RECT 598.235 -2.885 598.565 -2.555 ;
        RECT 596.875 -2.885 597.205 -2.555 ;
        RECT 595.515 -2.885 595.845 -2.555 ;
        RECT 594.155 -2.885 594.485 -2.555 ;
        RECT 592.795 -2.885 593.125 -2.555 ;
        RECT 591.435 -2.885 591.765 -2.555 ;
        RECT 590.075 -2.885 590.405 -2.555 ;
        RECT 588.715 -2.885 589.045 -2.555 ;
        RECT 587.355 -2.885 587.685 -2.555 ;
        RECT 585.995 -2.885 586.325 -2.555 ;
        RECT 584.635 -2.885 584.965 -2.555 ;
        RECT 583.275 -2.885 583.605 -2.555 ;
        RECT 581.915 -2.885 582.245 -2.555 ;
        RECT 580.555 -2.885 580.885 -2.555 ;
        RECT 579.195 -2.885 579.525 -2.555 ;
        RECT 577.835 -2.885 578.165 -2.555 ;
        RECT 576.475 -2.885 576.805 -2.555 ;
        RECT 575.115 -2.885 575.445 -2.555 ;
        RECT 573.755 -2.885 574.085 -2.555 ;
        RECT 572.395 -2.885 572.725 -2.555 ;
        RECT 571.035 -2.885 571.365 -2.555 ;
        RECT 569.675 -2.885 570.005 -2.555 ;
        RECT 568.315 -2.885 568.645 -2.555 ;
        RECT 566.955 -2.885 567.285 -2.555 ;
        RECT 565.595 -2.885 565.925 -2.555 ;
        RECT 564.235 -2.885 564.565 -2.555 ;
        RECT 562.875 -2.885 563.205 -2.555 ;
        RECT 561.515 -2.885 561.845 -2.555 ;
        RECT 560.155 -2.885 560.485 -2.555 ;
        RECT 558.795 -2.885 559.125 -2.555 ;
        RECT 557.435 -2.885 557.765 -2.555 ;
        RECT 556.075 -2.885 556.405 -2.555 ;
        RECT 554.715 -2.885 555.045 -2.555 ;
        RECT 553.355 -2.885 553.685 -2.555 ;
        RECT 551.995 -2.885 552.325 -2.555 ;
        RECT 550.635 -2.885 550.965 -2.555 ;
        RECT 549.275 -2.885 549.605 -2.555 ;
        RECT 547.915 -2.885 548.245 -2.555 ;
        RECT 546.555 -2.885 546.885 -2.555 ;
        RECT 545.195 -2.885 545.525 -2.555 ;
        RECT 543.835 -2.885 544.165 -2.555 ;
        RECT 542.475 -2.885 542.805 -2.555 ;
        RECT 541.115 -2.885 541.445 -2.555 ;
        RECT 539.755 -2.885 540.085 -2.555 ;
        RECT 538.395 -2.885 538.725 -2.555 ;
        RECT 537.035 -2.885 537.365 -2.555 ;
        RECT 535.675 -2.885 536.005 -2.555 ;
        RECT 534.315 -2.885 534.645 -2.555 ;
        RECT 532.955 -2.885 533.285 -2.555 ;
        RECT 531.595 -2.885 531.925 -2.555 ;
        RECT 530.235 -2.885 530.565 -2.555 ;
        RECT 528.875 -2.885 529.205 -2.555 ;
        RECT 527.515 -2.885 527.845 -2.555 ;
        RECT 526.155 -2.885 526.485 -2.555 ;
        RECT 524.795 -2.885 525.125 -2.555 ;
        RECT 523.435 -2.885 523.765 -2.555 ;
        RECT 522.075 -2.885 522.405 -2.555 ;
        RECT 520.715 -2.885 521.045 -2.555 ;
        RECT 519.355 -2.885 519.685 -2.555 ;
        RECT 517.995 -2.885 518.325 -2.555 ;
        RECT 516.635 -2.885 516.965 -2.555 ;
        RECT 515.275 -2.885 515.605 -2.555 ;
        RECT 513.915 -2.885 514.245 -2.555 ;
        RECT 512.555 -2.885 512.885 -2.555 ;
        RECT 511.195 -2.885 511.525 -2.555 ;
        RECT 509.835 -2.885 510.165 -2.555 ;
        RECT 508.475 -2.885 508.805 -2.555 ;
        RECT 507.115 -2.885 507.445 -2.555 ;
        RECT 505.755 -2.885 506.085 -2.555 ;
        RECT 504.395 -2.885 504.725 -2.555 ;
        RECT 503.035 -2.885 503.365 -2.555 ;
        RECT 501.675 -2.885 502.005 -2.555 ;
        RECT 500.315 -2.885 500.645 -2.555 ;
        RECT 498.955 -2.885 499.285 -2.555 ;
        RECT 497.595 -2.885 497.925 -2.555 ;
        RECT 496.235 -2.885 496.565 -2.555 ;
        RECT 494.875 -2.885 495.205 -2.555 ;
        RECT 493.515 -2.885 493.845 -2.555 ;
        RECT 492.155 -2.885 492.485 -2.555 ;
        RECT 490.795 -2.885 491.125 -2.555 ;
        RECT 489.435 -2.885 489.765 -2.555 ;
        RECT 488.075 -2.885 488.405 -2.555 ;
        RECT 486.715 -2.885 487.045 -2.555 ;
        RECT 485.355 -2.885 485.685 -2.555 ;
        RECT 483.995 -2.885 484.325 -2.555 ;
        RECT 482.635 -2.885 482.965 -2.555 ;
        RECT 481.275 -2.885 481.605 -2.555 ;
        RECT 479.915 -2.885 480.245 -2.555 ;
        RECT 478.555 -2.885 478.885 -2.555 ;
        RECT 477.195 -2.885 477.525 -2.555 ;
        RECT 475.835 -2.885 476.165 -2.555 ;
        RECT 474.475 -2.885 474.805 -2.555 ;
        RECT 473.115 -2.885 473.445 -2.555 ;
        RECT 471.755 -2.885 472.085 -2.555 ;
        RECT 470.395 -2.885 470.725 -2.555 ;
        RECT 469.035 -2.885 469.365 -2.555 ;
        RECT 467.675 -2.885 468.005 -2.555 ;
        RECT 466.315 -2.885 466.645 -2.555 ;
        RECT 464.955 -2.885 465.285 -2.555 ;
        RECT 463.595 -2.885 463.925 -2.555 ;
        RECT 462.235 -2.885 462.565 -2.555 ;
        RECT 460.875 -2.885 461.205 -2.555 ;
        RECT 459.515 -2.885 459.845 -2.555 ;
        RECT 458.155 -2.885 458.485 -2.555 ;
        RECT 456.795 -2.885 457.125 -2.555 ;
        RECT 455.435 -2.885 455.765 -2.555 ;
        RECT 454.075 -2.885 454.405 -2.555 ;
        RECT 452.715 -2.885 453.045 -2.555 ;
        RECT 451.355 -2.885 451.685 -2.555 ;
        RECT 449.995 -2.885 450.325 -2.555 ;
        RECT 448.635 -2.885 448.965 -2.555 ;
        RECT 447.275 -2.885 447.605 -2.555 ;
        RECT 445.915 -2.885 446.245 -2.555 ;
        RECT 444.555 -2.885 444.885 -2.555 ;
        RECT 443.195 -2.885 443.525 -2.555 ;
        RECT 441.835 -2.885 442.165 -2.555 ;
        RECT 440.475 -2.885 440.805 -2.555 ;
        RECT 439.115 -2.885 439.445 -2.555 ;
        RECT 437.755 -2.885 438.085 -2.555 ;
        RECT 436.395 -2.885 436.725 -2.555 ;
        RECT 435.035 -2.885 435.365 -2.555 ;
        RECT 433.675 -2.885 434.005 -2.555 ;
        RECT 432.315 -2.885 432.645 -2.555 ;
        RECT 430.955 -2.885 431.285 -2.555 ;
        RECT 429.595 -2.885 429.925 -2.555 ;
        RECT 428.235 -2.885 428.565 -2.555 ;
        RECT 426.875 -2.885 427.205 -2.555 ;
        RECT 425.515 -2.885 425.845 -2.555 ;
        RECT 424.155 -2.885 424.485 -2.555 ;
        RECT 422.795 -2.885 423.125 -2.555 ;
        RECT 421.435 -2.885 421.765 -2.555 ;
        RECT 420.075 -2.885 420.405 -2.555 ;
        RECT 418.715 -2.885 419.045 -2.555 ;
        RECT 417.355 -2.885 417.685 -2.555 ;
        RECT 415.995 -2.885 416.325 -2.555 ;
        RECT 414.635 -2.885 414.965 -2.555 ;
        RECT 413.275 -2.885 413.605 -2.555 ;
        RECT 411.915 -2.885 412.245 -2.555 ;
        RECT 410.555 -2.885 410.885 -2.555 ;
        RECT 409.195 -2.885 409.525 -2.555 ;
        RECT 407.835 -2.885 408.165 -2.555 ;
        RECT 406.475 -2.885 406.805 -2.555 ;
        RECT 405.115 -2.885 405.445 -2.555 ;
        RECT 403.755 -2.885 404.085 -2.555 ;
        RECT 402.395 -2.885 402.725 -2.555 ;
        RECT 401.035 -2.885 401.365 -2.555 ;
        RECT 399.675 -2.885 400.005 -2.555 ;
        RECT 398.315 -2.885 398.645 -2.555 ;
        RECT 396.955 -2.885 397.285 -2.555 ;
        RECT 395.595 -2.885 395.925 -2.555 ;
        RECT 394.235 -2.885 394.565 -2.555 ;
        RECT 392.875 -2.885 393.205 -2.555 ;
        RECT 391.515 -2.885 391.845 -2.555 ;
        RECT 390.155 -2.885 390.485 -2.555 ;
        RECT 388.795 -2.885 389.125 -2.555 ;
        RECT 387.435 -2.885 387.765 -2.555 ;
        RECT 386.075 -2.885 386.405 -2.555 ;
        RECT 384.715 -2.885 385.045 -2.555 ;
        RECT 383.355 -2.885 383.685 -2.555 ;
        RECT 381.995 -2.885 382.325 -2.555 ;
        RECT 380.635 -2.885 380.965 -2.555 ;
        RECT 379.275 -2.885 379.605 -2.555 ;
        RECT 377.915 -2.885 378.245 -2.555 ;
        RECT 376.555 -2.885 376.885 -2.555 ;
        RECT 375.195 -2.885 375.525 -2.555 ;
        RECT 373.835 -2.885 374.165 -2.555 ;
        RECT 372.475 -2.885 372.805 -2.555 ;
        RECT 371.115 -2.885 371.445 -2.555 ;
        RECT 369.755 -2.885 370.085 -2.555 ;
        RECT 368.395 -2.885 368.725 -2.555 ;
        RECT 367.035 -2.885 367.365 -2.555 ;
        RECT 365.675 -2.885 366.005 -2.555 ;
        RECT 364.315 -2.885 364.645 -2.555 ;
        RECT 362.955 -2.885 363.285 -2.555 ;
        RECT 361.595 -2.885 361.925 -2.555 ;
        RECT 360.235 -2.885 360.565 -2.555 ;
        RECT 358.875 -2.885 359.205 -2.555 ;
        RECT 357.515 -2.885 357.845 -2.555 ;
        RECT 356.155 -2.885 356.485 -2.555 ;
        RECT 354.795 -2.885 355.125 -2.555 ;
        RECT 353.435 -2.885 353.765 -2.555 ;
        RECT 352.075 -2.885 352.405 -2.555 ;
        RECT 350.715 -2.885 351.045 -2.555 ;
        RECT 349.355 -2.885 349.685 -2.555 ;
        RECT 347.995 -2.885 348.325 -2.555 ;
        RECT 346.635 -2.885 346.965 -2.555 ;
        RECT 345.275 -2.885 345.605 -2.555 ;
        RECT 343.915 -2.885 344.245 -2.555 ;
        RECT 342.555 -2.885 342.885 -2.555 ;
        RECT 341.195 -2.885 341.525 -2.555 ;
        RECT 339.835 -2.885 340.165 -2.555 ;
        RECT 338.475 -2.885 338.805 -2.555 ;
        RECT 337.115 -2.885 337.445 -2.555 ;
        RECT 335.755 -2.885 336.085 -2.555 ;
        RECT 334.395 -2.885 334.725 -2.555 ;
        RECT 333.035 -2.885 333.365 -2.555 ;
        RECT 331.675 -2.885 332.005 -2.555 ;
        RECT 330.315 -2.885 330.645 -2.555 ;
        RECT 328.955 -2.885 329.285 -2.555 ;
        RECT 327.595 -2.885 327.925 -2.555 ;
        RECT 326.235 -2.885 326.565 -2.555 ;
        RECT 324.875 -2.885 325.205 -2.555 ;
        RECT 323.515 -2.885 323.845 -2.555 ;
        RECT 322.155 -2.885 322.485 -2.555 ;
        RECT 320.795 -2.885 321.125 -2.555 ;
        RECT 319.435 -2.885 319.765 -2.555 ;
        RECT 318.075 -2.885 318.405 -2.555 ;
        RECT 316.715 -2.885 317.045 -2.555 ;
        RECT 315.355 -2.885 315.685 -2.555 ;
        RECT 313.995 -2.885 314.325 -2.555 ;
        RECT 312.635 -2.885 312.965 -2.555 ;
        RECT 311.275 -2.885 311.605 -2.555 ;
        RECT 309.915 -2.885 310.245 -2.555 ;
        RECT 308.555 -2.885 308.885 -2.555 ;
        RECT 307.195 -2.885 307.525 -2.555 ;
        RECT 305.835 -2.885 306.165 -2.555 ;
        RECT 304.475 -2.885 304.805 -2.555 ;
        RECT 303.115 -2.885 303.445 -2.555 ;
        RECT 301.755 -2.885 302.085 -2.555 ;
        RECT 300.395 -2.885 300.725 -2.555 ;
        RECT 299.035 -2.885 299.365 -2.555 ;
        RECT 297.675 -2.885 298.005 -2.555 ;
        RECT 296.315 -2.885 296.645 -2.555 ;
        RECT 294.955 -2.885 295.285 -2.555 ;
        RECT 293.595 -2.885 293.925 -2.555 ;
        RECT 292.235 -2.885 292.565 -2.555 ;
        RECT 290.875 -2.885 291.205 -2.555 ;
        RECT 289.515 -2.885 289.845 -2.555 ;
        RECT 288.155 -2.885 288.485 -2.555 ;
        RECT 286.795 -2.885 287.125 -2.555 ;
        RECT 285.435 -2.885 285.765 -2.555 ;
        RECT 284.075 -2.885 284.405 -2.555 ;
        RECT 282.715 -2.885 283.045 -2.555 ;
        RECT 281.355 -2.885 281.685 -2.555 ;
        RECT 279.995 -2.885 280.325 -2.555 ;
        RECT 278.635 -2.885 278.965 -2.555 ;
        RECT 277.275 -2.885 277.605 -2.555 ;
        RECT 275.915 -2.885 276.245 -2.555 ;
        RECT 274.555 -2.885 274.885 -2.555 ;
        RECT 273.195 -2.885 273.525 -2.555 ;
        RECT 271.835 -2.885 272.165 -2.555 ;
        RECT 270.475 -2.885 270.805 -2.555 ;
        RECT 269.115 -2.885 269.445 -2.555 ;
        RECT 267.755 -2.885 268.085 -2.555 ;
        RECT 266.395 -2.885 266.725 -2.555 ;
        RECT 265.035 -2.885 265.365 -2.555 ;
        RECT 263.675 -2.885 264.005 -2.555 ;
        RECT 262.315 -2.885 262.645 -2.555 ;
        RECT 260.955 -2.885 261.285 -2.555 ;
        RECT 259.595 -2.885 259.925 -2.555 ;
        RECT 258.235 -2.885 258.565 -2.555 ;
        RECT 256.875 -2.885 257.205 -2.555 ;
        RECT 255.515 -2.885 255.845 -2.555 ;
        RECT 254.155 -2.885 254.485 -2.555 ;
        RECT 252.795 -2.885 253.125 -2.555 ;
        RECT 251.435 -2.885 251.765 -2.555 ;
        RECT 250.075 -2.885 250.405 -2.555 ;
        RECT 248.715 -2.885 249.045 -2.555 ;
        RECT 247.355 -2.885 247.685 -2.555 ;
        RECT 245.995 -2.885 246.325 -2.555 ;
        RECT 244.635 -2.885 244.965 -2.555 ;
        RECT 243.275 -2.885 243.605 -2.555 ;
        RECT 241.915 -2.885 242.245 -2.555 ;
        RECT 240.555 -2.885 240.885 -2.555 ;
        RECT 239.195 -2.885 239.525 -2.555 ;
        RECT 237.835 -2.885 238.165 -2.555 ;
        RECT 236.475 -2.885 236.805 -2.555 ;
        RECT 235.115 -2.885 235.445 -2.555 ;
        RECT 233.755 -2.885 234.085 -2.555 ;
        RECT 232.395 -2.885 232.725 -2.555 ;
        RECT 231.035 -2.885 231.365 -2.555 ;
        RECT 229.675 -2.885 230.005 -2.555 ;
        RECT 228.315 -2.885 228.645 -2.555 ;
        RECT 226.955 -2.885 227.285 -2.555 ;
        RECT 225.595 -2.885 225.925 -2.555 ;
        RECT 224.235 -2.885 224.565 -2.555 ;
        RECT 222.875 -2.885 223.205 -2.555 ;
        RECT 221.515 -2.885 221.845 -2.555 ;
        RECT 220.155 -2.885 220.485 -2.555 ;
        RECT 218.795 -2.885 219.125 -2.555 ;
        RECT 217.435 -2.885 217.765 -2.555 ;
        RECT 216.075 -2.885 216.405 -2.555 ;
        RECT 214.715 -2.885 215.045 -2.555 ;
        RECT 213.355 -2.885 213.685 -2.555 ;
        RECT 211.995 -2.885 212.325 -2.555 ;
        RECT 210.635 -2.885 210.965 -2.555 ;
        RECT 209.275 -2.885 209.605 -2.555 ;
        RECT 207.915 -2.885 208.245 -2.555 ;
        RECT 206.555 -2.885 206.885 -2.555 ;
        RECT 205.195 -2.885 205.525 -2.555 ;
        RECT 203.835 -2.885 204.165 -2.555 ;
        RECT 202.475 -2.885 202.805 -2.555 ;
        RECT 201.115 -2.885 201.445 -2.555 ;
        RECT 199.755 -2.885 200.085 -2.555 ;
        RECT 198.395 -2.885 198.725 -2.555 ;
        RECT 197.035 -2.885 197.365 -2.555 ;
        RECT 195.675 -2.885 196.005 -2.555 ;
        RECT 194.315 -2.885 194.645 -2.555 ;
        RECT 192.955 -2.885 193.285 -2.555 ;
        RECT 191.595 -2.885 191.925 -2.555 ;
        RECT 190.235 -2.885 190.565 -2.555 ;
        RECT 188.875 -2.885 189.205 -2.555 ;
        RECT 187.515 -2.885 187.845 -2.555 ;
        RECT 186.155 -2.885 186.485 -2.555 ;
        RECT 184.795 -2.885 185.125 -2.555 ;
        RECT 183.435 -2.885 183.765 -2.555 ;
        RECT 182.075 -2.885 182.405 -2.555 ;
        RECT 180.715 -2.885 181.045 -2.555 ;
        RECT 179.355 -2.885 179.685 -2.555 ;
        RECT 177.995 -2.885 178.325 -2.555 ;
        RECT 176.635 -2.885 176.965 -2.555 ;
        RECT 175.275 -2.885 175.605 -2.555 ;
        RECT 173.915 -2.885 174.245 -2.555 ;
        RECT 172.555 -2.885 172.885 -2.555 ;
        RECT 171.195 -2.885 171.525 -2.555 ;
        RECT 169.835 -2.885 170.165 -2.555 ;
        RECT 168.475 -2.885 168.805 -2.555 ;
        RECT 167.115 -2.885 167.445 -2.555 ;
        RECT 165.755 -2.885 166.085 -2.555 ;
        RECT 164.395 -2.885 164.725 -2.555 ;
        RECT 163.035 -2.885 163.365 -2.555 ;
        RECT 161.675 -2.885 162.005 -2.555 ;
        RECT 160.315 -2.885 160.645 -2.555 ;
        RECT 158.955 -2.885 159.285 -2.555 ;
        RECT 157.595 -2.885 157.925 -2.555 ;
        RECT 156.235 -2.885 156.565 -2.555 ;
        RECT 154.875 -2.885 155.205 -2.555 ;
        RECT 153.515 -2.885 153.845 -2.555 ;
        RECT 152.155 -2.885 152.485 -2.555 ;
        RECT 150.795 -2.885 151.125 -2.555 ;
        RECT 149.435 -2.885 149.765 -2.555 ;
        RECT 148.075 -2.885 148.405 -2.555 ;
        RECT 146.715 -2.885 147.045 -2.555 ;
        RECT 145.355 -2.885 145.685 -2.555 ;
        RECT 143.995 -2.885 144.325 -2.555 ;
        RECT 142.635 -2.885 142.965 -2.555 ;
        RECT 141.275 -2.885 141.605 -2.555 ;
        RECT 139.915 -2.885 140.245 -2.555 ;
        RECT 138.555 -2.885 138.885 -2.555 ;
        RECT 137.195 -2.885 137.525 -2.555 ;
        RECT 135.835 -2.885 136.165 -2.555 ;
        RECT 134.475 -2.885 134.805 -2.555 ;
        RECT 133.115 -2.885 133.445 -2.555 ;
        RECT 131.755 -2.885 132.085 -2.555 ;
        RECT 130.395 -2.885 130.725 -2.555 ;
        RECT 129.035 -2.885 129.365 -2.555 ;
        RECT 127.675 -2.885 128.005 -2.555 ;
        RECT 126.315 -2.885 126.645 -2.555 ;
        RECT 124.955 -2.885 125.285 -2.555 ;
        RECT 123.595 -2.885 123.925 -2.555 ;
        RECT 122.235 -2.885 122.565 -2.555 ;
        RECT 120.875 -2.885 121.205 -2.555 ;
        RECT 119.515 -2.885 119.845 -2.555 ;
        RECT 118.155 -2.885 118.485 -2.555 ;
        RECT 116.795 -2.885 117.125 -2.555 ;
        RECT 115.435 -2.885 115.765 -2.555 ;
        RECT 114.075 -2.885 114.405 -2.555 ;
        RECT 112.715 -2.885 113.045 -2.555 ;
        RECT 111.355 -2.885 111.685 -2.555 ;
        RECT 109.995 -2.885 110.325 -2.555 ;
        RECT 108.635 -2.885 108.965 -2.555 ;
        RECT 107.275 -2.885 107.605 -2.555 ;
        RECT 105.915 -2.885 106.245 -2.555 ;
        RECT 104.555 -2.885 104.885 -2.555 ;
        RECT 103.195 -2.885 103.525 -2.555 ;
        RECT 101.835 -2.885 102.165 -2.555 ;
        RECT 100.475 -2.885 100.805 -2.555 ;
        RECT 99.115 -2.885 99.445 -2.555 ;
        RECT 97.755 -2.885 98.085 -2.555 ;
        RECT 96.395 -2.885 96.725 -2.555 ;
        RECT 95.035 -2.885 95.365 -2.555 ;
        RECT 93.675 -2.885 94.005 -2.555 ;
        RECT 92.315 -2.885 92.645 -2.555 ;
        RECT 90.955 -2.885 91.285 -2.555 ;
        RECT 89.595 -2.885 89.925 -2.555 ;
        RECT 88.235 -2.885 88.565 -2.555 ;
        RECT 86.875 -2.885 87.205 -2.555 ;
        RECT 85.515 -2.885 85.845 -2.555 ;
        RECT 84.155 -2.885 84.485 -2.555 ;
        RECT 82.795 -2.885 83.125 -2.555 ;
        RECT 81.435 -2.885 81.765 -2.555 ;
        RECT 80.075 -2.885 80.405 -2.555 ;
        RECT 78.715 -2.885 79.045 -2.555 ;
        RECT 77.355 -2.885 77.685 -2.555 ;
        RECT 75.995 -2.885 76.325 -2.555 ;
        RECT 74.635 -2.885 74.965 -2.555 ;
        RECT 73.275 -2.885 73.605 -2.555 ;
        RECT 71.915 -2.885 72.245 -2.555 ;
        RECT 70.555 -2.885 70.885 -2.555 ;
        RECT 69.195 -2.885 69.525 -2.555 ;
        RECT 67.835 -2.885 68.165 -2.555 ;
        RECT 66.475 -2.885 66.805 -2.555 ;
        RECT 65.115 -2.885 65.445 -2.555 ;
        RECT 63.755 -2.885 64.085 -2.555 ;
        RECT 62.395 -2.885 62.725 -2.555 ;
        RECT 61.035 -2.885 61.365 -2.555 ;
        RECT 59.675 -2.885 60.005 -2.555 ;
        RECT 58.315 -2.885 58.645 -2.555 ;
        RECT 56.955 -2.885 57.285 -2.555 ;
        RECT 55.595 -2.885 55.925 -2.555 ;
        RECT 54.235 -2.885 54.565 -2.555 ;
        RECT 52.875 -2.885 53.205 -2.555 ;
        RECT 51.515 -2.885 51.845 -2.555 ;
        RECT 50.155 -2.885 50.485 -2.555 ;
        RECT 48.795 -2.885 49.125 -2.555 ;
        RECT 47.435 -2.885 47.765 -2.555 ;
        RECT 46.075 -2.885 46.405 -2.555 ;
        RECT 44.715 -2.885 45.045 -2.555 ;
        RECT 43.355 -2.885 43.685 -2.555 ;
        RECT 41.995 -2.885 42.325 -2.555 ;
        RECT 40.635 -2.885 40.965 -2.555 ;
        RECT 39.275 -2.885 39.605 -2.555 ;
        RECT 37.915 -2.885 38.245 -2.555 ;
        RECT 36.555 -2.885 36.885 -2.555 ;
        RECT 35.195 -2.885 35.525 -2.555 ;
        RECT 33.835 -2.885 34.165 -2.555 ;
        RECT 32.475 -2.885 32.805 -2.555 ;
        RECT 31.115 -2.885 31.445 -2.555 ;
        RECT 29.755 -2.885 30.085 -2.555 ;
        RECT 28.395 -2.885 28.725 -2.555 ;
        RECT 27.035 -2.885 27.365 -2.555 ;
        RECT 25.675 -2.885 26.005 -2.555 ;
        RECT 24.315 -2.885 24.645 -2.555 ;
        RECT 22.955 -2.885 23.285 -2.555 ;
        RECT 21.595 -2.885 21.925 -2.555 ;
        RECT 20.235 -2.885 20.565 -2.555 ;
        RECT 18.875 -2.885 19.205 -2.555 ;
        RECT 17.515 -2.885 17.845 -2.555 ;
        RECT 16.155 -2.885 16.485 -2.555 ;
        RECT 14.795 -2.885 15.125 -2.555 ;
        RECT 13.435 -2.885 13.765 -2.555 ;
        RECT 12.075 -2.885 12.405 -2.555 ;
        RECT 10.715 -2.885 11.045 -2.555 ;
        RECT 9.355 -2.885 9.685 -2.555 ;
        RECT 7.995 -2.885 8.325 -2.555 ;
        RECT 6.635 -2.885 6.965 -2.555 ;
        RECT 5.275 -2.885 5.605 -2.555 ;
        RECT 3.915 -2.885 4.245 -2.555 ;
        RECT 2.555 -2.885 2.885 -2.555 ;
        RECT 1.195 -2.885 1.525 -2.555 ;
        RECT -0.165 -2.885 0.165 -2.555 ;
        RECT -1.525 -2.885 -1.195 -2.555 ;
        RECT -1.525 -2.88 678.475 -2.56 ;
        RECT 677.115 -2.885 677.445 -2.555 ;
        RECT 675.755 -2.885 676.085 -2.555 ;
        RECT 674.395 -2.885 674.725 -2.555 ;
        RECT 673.035 -2.885 673.365 -2.555 ;
        RECT 671.675 -2.885 672.005 -2.555 ;
        RECT 670.315 -2.885 670.645 -2.555 ;
        RECT 668.955 -2.885 669.285 -2.555 ;
        RECT 667.595 -2.885 667.925 -2.555 ;
        RECT 666.235 -2.885 666.565 -2.555 ;
        RECT 664.875 -2.885 665.205 -2.555 ;
        RECT 663.515 -2.885 663.845 -2.555 ;
        RECT 662.155 -2.885 662.485 -2.555 ;
        RECT 660.795 -2.885 661.125 -2.555 ;
        RECT 659.435 -2.885 659.765 -2.555 ;
        RECT 658.075 -2.885 658.405 -2.555 ;
        RECT 954.555 -2.885 954.885 -2.555 ;
        RECT 678.475 -2.88 954.885 -2.56 ;
        RECT 953.195 -2.885 953.525 -2.555 ;
        RECT 951.835 -2.885 952.165 -2.555 ;
        RECT 950.475 -2.885 950.805 -2.555 ;
        RECT 949.115 -2.885 949.445 -2.555 ;
        RECT 947.755 -2.885 948.085 -2.555 ;
        RECT 946.395 -2.885 946.725 -2.555 ;
        RECT 945.035 -2.885 945.365 -2.555 ;
        RECT 943.675 -2.885 944.005 -2.555 ;
        RECT 942.315 -2.885 942.645 -2.555 ;
        RECT 940.955 -2.885 941.285 -2.555 ;
        RECT 939.595 -2.885 939.925 -2.555 ;
        RECT 938.235 -2.885 938.565 -2.555 ;
        RECT 936.875 -2.885 937.205 -2.555 ;
        RECT 935.515 -2.885 935.845 -2.555 ;
        RECT 934.155 -2.885 934.485 -2.555 ;
        RECT 932.795 -2.885 933.125 -2.555 ;
        RECT 931.435 -2.885 931.765 -2.555 ;
        RECT 930.075 -2.885 930.405 -2.555 ;
        RECT 928.715 -2.885 929.045 -2.555 ;
        RECT 927.355 -2.885 927.685 -2.555 ;
        RECT 925.995 -2.885 926.325 -2.555 ;
        RECT 924.635 -2.885 924.965 -2.555 ;
        RECT 923.275 -2.885 923.605 -2.555 ;
        RECT 921.915 -2.885 922.245 -2.555 ;
        RECT 920.555 -2.885 920.885 -2.555 ;
        RECT 919.195 -2.885 919.525 -2.555 ;
        RECT 917.835 -2.885 918.165 -2.555 ;
        RECT 916.475 -2.885 916.805 -2.555 ;
        RECT 915.115 -2.885 915.445 -2.555 ;
        RECT 913.755 -2.885 914.085 -2.555 ;
        RECT 912.395 -2.885 912.725 -2.555 ;
        RECT 911.035 -2.885 911.365 -2.555 ;
        RECT 909.675 -2.885 910.005 -2.555 ;
        RECT 908.315 -2.885 908.645 -2.555 ;
        RECT 906.955 -2.885 907.285 -2.555 ;
        RECT 905.595 -2.885 905.925 -2.555 ;
        RECT 904.235 -2.885 904.565 -2.555 ;
        RECT 902.875 -2.885 903.205 -2.555 ;
        RECT 901.515 -2.885 901.845 -2.555 ;
        RECT 900.155 -2.885 900.485 -2.555 ;
        RECT 898.795 -2.885 899.125 -2.555 ;
        RECT 897.435 -2.885 897.765 -2.555 ;
        RECT 896.075 -2.885 896.405 -2.555 ;
        RECT 894.715 -2.885 895.045 -2.555 ;
        RECT 893.355 -2.885 893.685 -2.555 ;
        RECT 891.995 -2.885 892.325 -2.555 ;
        RECT 890.635 -2.885 890.965 -2.555 ;
        RECT 889.275 -2.885 889.605 -2.555 ;
        RECT 887.915 -2.885 888.245 -2.555 ;
        RECT 886.555 -2.885 886.885 -2.555 ;
        RECT 885.195 -2.885 885.525 -2.555 ;
        RECT 883.835 -2.885 884.165 -2.555 ;
        RECT 882.475 -2.885 882.805 -2.555 ;
        RECT 881.115 -2.885 881.445 -2.555 ;
        RECT 879.755 -2.885 880.085 -2.555 ;
        RECT 878.395 -2.885 878.725 -2.555 ;
        RECT 877.035 -2.885 877.365 -2.555 ;
        RECT 875.675 -2.885 876.005 -2.555 ;
        RECT 874.315 -2.885 874.645 -2.555 ;
        RECT 872.955 -2.885 873.285 -2.555 ;
        RECT 871.595 -2.885 871.925 -2.555 ;
        RECT 870.235 -2.885 870.565 -2.555 ;
        RECT 868.875 -2.885 869.205 -2.555 ;
        RECT 867.515 -2.885 867.845 -2.555 ;
        RECT 866.155 -2.885 866.485 -2.555 ;
        RECT 864.795 -2.885 865.125 -2.555 ;
        RECT 863.435 -2.885 863.765 -2.555 ;
        RECT 862.075 -2.885 862.405 -2.555 ;
        RECT 860.715 -2.885 861.045 -2.555 ;
        RECT 859.355 -2.885 859.685 -2.555 ;
        RECT 857.995 -2.885 858.325 -2.555 ;
        RECT 856.635 -2.885 856.965 -2.555 ;
        RECT 855.275 -2.885 855.605 -2.555 ;
        RECT 853.915 -2.885 854.245 -2.555 ;
        RECT 852.555 -2.885 852.885 -2.555 ;
        RECT 851.195 -2.885 851.525 -2.555 ;
        RECT 849.835 -2.885 850.165 -2.555 ;
        RECT 848.475 -2.885 848.805 -2.555 ;
        RECT 847.115 -2.885 847.445 -2.555 ;
        RECT 845.755 -2.885 846.085 -2.555 ;
        RECT 844.395 -2.885 844.725 -2.555 ;
        RECT 843.035 -2.885 843.365 -2.555 ;
        RECT 841.675 -2.885 842.005 -2.555 ;
        RECT 840.315 -2.885 840.645 -2.555 ;
        RECT 838.955 -2.885 839.285 -2.555 ;
        RECT 837.595 -2.885 837.925 -2.555 ;
        RECT 836.235 -2.885 836.565 -2.555 ;
        RECT 834.875 -2.885 835.205 -2.555 ;
        RECT 833.515 -2.885 833.845 -2.555 ;
        RECT 832.155 -2.885 832.485 -2.555 ;
        RECT 830.795 -2.885 831.125 -2.555 ;
        RECT 829.435 -2.885 829.765 -2.555 ;
        RECT 828.075 -2.885 828.405 -2.555 ;
        RECT 826.715 -2.885 827.045 -2.555 ;
        RECT 825.355 -2.885 825.685 -2.555 ;
        RECT 823.995 -2.885 824.325 -2.555 ;
        RECT 822.635 -2.885 822.965 -2.555 ;
        RECT 821.275 -2.885 821.605 -2.555 ;
        RECT 819.915 -2.885 820.245 -2.555 ;
        RECT 818.555 -2.885 818.885 -2.555 ;
        RECT 817.195 -2.885 817.525 -2.555 ;
        RECT 815.835 -2.885 816.165 -2.555 ;
        RECT 814.475 -2.885 814.805 -2.555 ;
        RECT 813.115 -2.885 813.445 -2.555 ;
        RECT 811.755 -2.885 812.085 -2.555 ;
        RECT 810.395 -2.885 810.725 -2.555 ;
        RECT 809.035 -2.885 809.365 -2.555 ;
        RECT 807.675 -2.885 808.005 -2.555 ;
        RECT 806.315 -2.885 806.645 -2.555 ;
        RECT 804.955 -2.885 805.285 -2.555 ;
        RECT 803.595 -2.885 803.925 -2.555 ;
        RECT 802.235 -2.885 802.565 -2.555 ;
        RECT 800.875 -2.885 801.205 -2.555 ;
        RECT 799.515 -2.885 799.845 -2.555 ;
        RECT 798.155 -2.885 798.485 -2.555 ;
        RECT 796.795 -2.885 797.125 -2.555 ;
        RECT 795.435 -2.885 795.765 -2.555 ;
        RECT 794.075 -2.885 794.405 -2.555 ;
        RECT 792.715 -2.885 793.045 -2.555 ;
        RECT 791.355 -2.885 791.685 -2.555 ;
        RECT 789.995 -2.885 790.325 -2.555 ;
        RECT 788.635 -2.885 788.965 -2.555 ;
        RECT 787.275 -2.885 787.605 -2.555 ;
        RECT 785.915 -2.885 786.245 -2.555 ;
        RECT 784.555 -2.885 784.885 -2.555 ;
        RECT 783.195 -2.885 783.525 -2.555 ;
        RECT 781.835 -2.885 782.165 -2.555 ;
        RECT 780.475 -2.885 780.805 -2.555 ;
        RECT 779.115 -2.885 779.445 -2.555 ;
        RECT 777.755 -2.885 778.085 -2.555 ;
        RECT 776.395 -2.885 776.725 -2.555 ;
        RECT 775.035 -2.885 775.365 -2.555 ;
        RECT 773.675 -2.885 774.005 -2.555 ;
        RECT 772.315 -2.885 772.645 -2.555 ;
        RECT 770.955 -2.885 771.285 -2.555 ;
        RECT 769.595 -2.885 769.925 -2.555 ;
        RECT 768.235 -2.885 768.565 -2.555 ;
        RECT 766.875 -2.885 767.205 -2.555 ;
        RECT 765.515 -2.885 765.845 -2.555 ;
        RECT 764.155 -2.885 764.485 -2.555 ;
        RECT 762.795 -2.885 763.125 -2.555 ;
        RECT 761.435 -2.885 761.765 -2.555 ;
        RECT 760.075 -2.885 760.405 -2.555 ;
        RECT 758.715 -2.885 759.045 -2.555 ;
        RECT 757.355 -2.885 757.685 -2.555 ;
        RECT 755.995 -2.885 756.325 -2.555 ;
        RECT 754.635 -2.885 754.965 -2.555 ;
        RECT 753.275 -2.885 753.605 -2.555 ;
        RECT 751.915 -2.885 752.245 -2.555 ;
        RECT 750.555 -2.885 750.885 -2.555 ;
        RECT 749.195 -2.885 749.525 -2.555 ;
        RECT 747.835 -2.885 748.165 -2.555 ;
        RECT 746.475 -2.885 746.805 -2.555 ;
        RECT 745.115 -2.885 745.445 -2.555 ;
        RECT 743.755 -2.885 744.085 -2.555 ;
        RECT 742.395 -2.885 742.725 -2.555 ;
        RECT 741.035 -2.885 741.365 -2.555 ;
        RECT 739.675 -2.885 740.005 -2.555 ;
        RECT 738.315 -2.885 738.645 -2.555 ;
        RECT 736.955 -2.885 737.285 -2.555 ;
        RECT 735.595 -2.885 735.925 -2.555 ;
        RECT 734.235 -2.885 734.565 -2.555 ;
        RECT 732.875 -2.885 733.205 -2.555 ;
        RECT 731.515 -2.885 731.845 -2.555 ;
        RECT 730.155 -2.885 730.485 -2.555 ;
        RECT 728.795 -2.885 729.125 -2.555 ;
        RECT 727.435 -2.885 727.765 -2.555 ;
        RECT 726.075 -2.885 726.405 -2.555 ;
        RECT 724.715 -2.885 725.045 -2.555 ;
        RECT 723.355 -2.885 723.685 -2.555 ;
        RECT 721.995 -2.885 722.325 -2.555 ;
        RECT 720.635 -2.885 720.965 -2.555 ;
        RECT 719.275 -2.885 719.605 -2.555 ;
        RECT 717.915 -2.885 718.245 -2.555 ;
        RECT 716.555 -2.885 716.885 -2.555 ;
        RECT 715.195 -2.885 715.525 -2.555 ;
        RECT 713.835 -2.885 714.165 -2.555 ;
        RECT 712.475 -2.885 712.805 -2.555 ;
        RECT 711.115 -2.885 711.445 -2.555 ;
        RECT 709.755 -2.885 710.085 -2.555 ;
        RECT 708.395 -2.885 708.725 -2.555 ;
        RECT 707.035 -2.885 707.365 -2.555 ;
        RECT 705.675 -2.885 706.005 -2.555 ;
        RECT 704.315 -2.885 704.645 -2.555 ;
        RECT 702.955 -2.885 703.285 -2.555 ;
        RECT 701.595 -2.885 701.925 -2.555 ;
        RECT 700.235 -2.885 700.565 -2.555 ;
        RECT 698.875 -2.885 699.205 -2.555 ;
        RECT 697.515 -2.885 697.845 -2.555 ;
        RECT 696.155 -2.885 696.485 -2.555 ;
        RECT 694.795 -2.885 695.125 -2.555 ;
        RECT 693.435 -2.885 693.765 -2.555 ;
        RECT 692.075 -2.885 692.405 -2.555 ;
        RECT 690.715 -2.885 691.045 -2.555 ;
        RECT 689.355 -2.885 689.685 -2.555 ;
        RECT 687.995 -2.885 688.325 -2.555 ;
        RECT 686.635 -2.885 686.965 -2.555 ;
        RECT 685.275 -2.885 685.605 -2.555 ;
        RECT 683.915 -2.885 684.245 -2.555 ;
        RECT 682.555 -2.885 682.885 -2.555 ;
        RECT 681.195 -2.885 681.525 -2.555 ;
        RECT 679.835 -2.885 680.165 -2.555 ;
        RECT 678.475 -2.885 678.805 -2.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.92 -26 677.44 -25.68 ;
        RECT 675.755 -26.005 676.085 -25.675 ;
        RECT 674.395 -26.005 674.725 -25.675 ;
        RECT 671.675 -26.005 672.005 -25.675 ;
        RECT 670.315 -26.005 670.645 -25.675 ;
        RECT 668.955 -26.005 669.285 -25.675 ;
        RECT 667.595 -26.005 667.925 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 1.2 678.475 1.52 ;
        RECT 677.115 1.195 677.445 1.525 ;
        RECT 675.755 1.195 676.085 1.525 ;
        RECT 674.395 1.195 674.725 1.525 ;
        RECT 673.035 1.195 673.365 1.525 ;
        RECT 671.675 1.195 672.005 1.525 ;
        RECT 670.315 1.195 670.645 1.525 ;
        RECT 668.955 1.195 669.285 1.525 ;
        RECT 667.595 1.195 667.925 1.525 ;
        RECT 666.235 1.195 666.565 1.525 ;
        RECT 664.875 1.195 665.205 1.525 ;
        RECT 663.515 1.195 663.845 1.525 ;
        RECT 662.155 1.195 662.485 1.525 ;
        RECT 660.795 1.195 661.125 1.525 ;
        RECT 659.435 1.195 659.765 1.525 ;
        RECT 658.075 1.195 658.405 1.525 ;
        RECT 656.715 1.195 657.045 1.525 ;
        RECT 655.355 1.195 655.685 1.525 ;
        RECT 653.995 1.195 654.325 1.525 ;
        RECT 652.635 1.195 652.965 1.525 ;
        RECT 651.275 1.195 651.605 1.525 ;
        RECT 649.915 1.195 650.245 1.525 ;
        RECT 648.555 1.195 648.885 1.525 ;
        RECT 647.195 1.195 647.525 1.525 ;
        RECT 645.835 1.195 646.165 1.525 ;
        RECT 644.475 1.195 644.805 1.525 ;
        RECT 643.115 1.195 643.445 1.525 ;
        RECT 641.755 1.195 642.085 1.525 ;
        RECT 640.395 1.195 640.725 1.525 ;
        RECT 639.035 1.195 639.365 1.525 ;
        RECT 637.675 1.195 638.005 1.525 ;
        RECT 636.315 1.195 636.645 1.525 ;
        RECT 634.955 1.195 635.285 1.525 ;
        RECT 633.595 1.195 633.925 1.525 ;
        RECT 632.235 1.195 632.565 1.525 ;
        RECT 630.875 1.195 631.205 1.525 ;
        RECT 629.515 1.195 629.845 1.525 ;
        RECT 628.155 1.195 628.485 1.525 ;
        RECT 626.795 1.195 627.125 1.525 ;
        RECT 625.435 1.195 625.765 1.525 ;
        RECT 624.075 1.195 624.405 1.525 ;
        RECT 622.715 1.195 623.045 1.525 ;
        RECT 621.355 1.195 621.685 1.525 ;
        RECT 619.995 1.195 620.325 1.525 ;
        RECT 618.635 1.195 618.965 1.525 ;
        RECT 617.275 1.195 617.605 1.525 ;
        RECT 615.915 1.195 616.245 1.525 ;
        RECT 614.555 1.195 614.885 1.525 ;
        RECT 613.195 1.195 613.525 1.525 ;
        RECT 611.835 1.195 612.165 1.525 ;
        RECT 610.475 1.195 610.805 1.525 ;
        RECT 609.115 1.195 609.445 1.525 ;
        RECT 607.755 1.195 608.085 1.525 ;
        RECT 606.395 1.195 606.725 1.525 ;
        RECT 605.035 1.195 605.365 1.525 ;
        RECT 603.675 1.195 604.005 1.525 ;
        RECT 602.315 1.195 602.645 1.525 ;
        RECT 600.955 1.195 601.285 1.525 ;
        RECT 599.595 1.195 599.925 1.525 ;
        RECT 598.235 1.195 598.565 1.525 ;
        RECT 596.875 1.195 597.205 1.525 ;
        RECT 595.515 1.195 595.845 1.525 ;
        RECT 594.155 1.195 594.485 1.525 ;
        RECT 592.795 1.195 593.125 1.525 ;
        RECT 591.435 1.195 591.765 1.525 ;
        RECT 590.075 1.195 590.405 1.525 ;
        RECT 588.715 1.195 589.045 1.525 ;
        RECT 587.355 1.195 587.685 1.525 ;
        RECT 585.995 1.195 586.325 1.525 ;
        RECT 584.635 1.195 584.965 1.525 ;
        RECT 583.275 1.195 583.605 1.525 ;
        RECT 581.915 1.195 582.245 1.525 ;
        RECT 580.555 1.195 580.885 1.525 ;
        RECT 579.195 1.195 579.525 1.525 ;
        RECT 577.835 1.195 578.165 1.525 ;
        RECT 576.475 1.195 576.805 1.525 ;
        RECT 575.115 1.195 575.445 1.525 ;
        RECT 573.755 1.195 574.085 1.525 ;
        RECT 572.395 1.195 572.725 1.525 ;
        RECT 571.035 1.195 571.365 1.525 ;
        RECT 569.675 1.195 570.005 1.525 ;
        RECT 568.315 1.195 568.645 1.525 ;
        RECT 566.955 1.195 567.285 1.525 ;
        RECT 565.595 1.195 565.925 1.525 ;
        RECT 564.235 1.195 564.565 1.525 ;
        RECT 562.875 1.195 563.205 1.525 ;
        RECT 561.515 1.195 561.845 1.525 ;
        RECT 560.155 1.195 560.485 1.525 ;
        RECT 558.795 1.195 559.125 1.525 ;
        RECT 557.435 1.195 557.765 1.525 ;
        RECT 556.075 1.195 556.405 1.525 ;
        RECT 554.715 1.195 555.045 1.525 ;
        RECT 553.355 1.195 553.685 1.525 ;
        RECT 551.995 1.195 552.325 1.525 ;
        RECT 550.635 1.195 550.965 1.525 ;
        RECT 549.275 1.195 549.605 1.525 ;
        RECT 547.915 1.195 548.245 1.525 ;
        RECT 546.555 1.195 546.885 1.525 ;
        RECT 545.195 1.195 545.525 1.525 ;
        RECT 543.835 1.195 544.165 1.525 ;
        RECT 542.475 1.195 542.805 1.525 ;
        RECT 541.115 1.195 541.445 1.525 ;
        RECT 539.755 1.195 540.085 1.525 ;
        RECT 538.395 1.195 538.725 1.525 ;
        RECT 537.035 1.195 537.365 1.525 ;
        RECT 535.675 1.195 536.005 1.525 ;
        RECT 534.315 1.195 534.645 1.525 ;
        RECT 532.955 1.195 533.285 1.525 ;
        RECT 531.595 1.195 531.925 1.525 ;
        RECT 530.235 1.195 530.565 1.525 ;
        RECT 528.875 1.195 529.205 1.525 ;
        RECT 527.515 1.195 527.845 1.525 ;
        RECT 526.155 1.195 526.485 1.525 ;
        RECT 524.795 1.195 525.125 1.525 ;
        RECT 523.435 1.195 523.765 1.525 ;
        RECT 522.075 1.195 522.405 1.525 ;
        RECT 520.715 1.195 521.045 1.525 ;
        RECT 519.355 1.195 519.685 1.525 ;
        RECT 517.995 1.195 518.325 1.525 ;
        RECT 516.635 1.195 516.965 1.525 ;
        RECT 515.275 1.195 515.605 1.525 ;
        RECT 513.915 1.195 514.245 1.525 ;
        RECT 512.555 1.195 512.885 1.525 ;
        RECT 511.195 1.195 511.525 1.525 ;
        RECT 509.835 1.195 510.165 1.525 ;
        RECT 508.475 1.195 508.805 1.525 ;
        RECT 507.115 1.195 507.445 1.525 ;
        RECT 505.755 1.195 506.085 1.525 ;
        RECT 504.395 1.195 504.725 1.525 ;
        RECT 503.035 1.195 503.365 1.525 ;
        RECT 501.675 1.195 502.005 1.525 ;
        RECT 500.315 1.195 500.645 1.525 ;
        RECT 498.955 1.195 499.285 1.525 ;
        RECT 497.595 1.195 497.925 1.525 ;
        RECT 496.235 1.195 496.565 1.525 ;
        RECT 494.875 1.195 495.205 1.525 ;
        RECT 493.515 1.195 493.845 1.525 ;
        RECT 492.155 1.195 492.485 1.525 ;
        RECT 490.795 1.195 491.125 1.525 ;
        RECT 489.435 1.195 489.765 1.525 ;
        RECT 488.075 1.195 488.405 1.525 ;
        RECT 486.715 1.195 487.045 1.525 ;
        RECT 485.355 1.195 485.685 1.525 ;
        RECT 483.995 1.195 484.325 1.525 ;
        RECT 482.635 1.195 482.965 1.525 ;
        RECT 481.275 1.195 481.605 1.525 ;
        RECT 479.915 1.195 480.245 1.525 ;
        RECT 478.555 1.195 478.885 1.525 ;
        RECT 477.195 1.195 477.525 1.525 ;
        RECT 475.835 1.195 476.165 1.525 ;
        RECT 474.475 1.195 474.805 1.525 ;
        RECT 473.115 1.195 473.445 1.525 ;
        RECT 471.755 1.195 472.085 1.525 ;
        RECT 470.395 1.195 470.725 1.525 ;
        RECT 469.035 1.195 469.365 1.525 ;
        RECT 467.675 1.195 468.005 1.525 ;
        RECT 466.315 1.195 466.645 1.525 ;
        RECT 464.955 1.195 465.285 1.525 ;
        RECT 463.595 1.195 463.925 1.525 ;
        RECT 462.235 1.195 462.565 1.525 ;
        RECT 460.875 1.195 461.205 1.525 ;
        RECT 459.515 1.195 459.845 1.525 ;
        RECT 458.155 1.195 458.485 1.525 ;
        RECT 456.795 1.195 457.125 1.525 ;
        RECT 455.435 1.195 455.765 1.525 ;
        RECT 454.075 1.195 454.405 1.525 ;
        RECT 452.715 1.195 453.045 1.525 ;
        RECT 451.355 1.195 451.685 1.525 ;
        RECT 449.995 1.195 450.325 1.525 ;
        RECT 448.635 1.195 448.965 1.525 ;
        RECT 447.275 1.195 447.605 1.525 ;
        RECT 445.915 1.195 446.245 1.525 ;
        RECT 444.555 1.195 444.885 1.525 ;
        RECT 443.195 1.195 443.525 1.525 ;
        RECT 441.835 1.195 442.165 1.525 ;
        RECT 440.475 1.195 440.805 1.525 ;
        RECT 439.115 1.195 439.445 1.525 ;
        RECT 437.755 1.195 438.085 1.525 ;
        RECT 436.395 1.195 436.725 1.525 ;
        RECT 435.035 1.195 435.365 1.525 ;
        RECT 433.675 1.195 434.005 1.525 ;
        RECT 432.315 1.195 432.645 1.525 ;
        RECT 430.955 1.195 431.285 1.525 ;
        RECT 429.595 1.195 429.925 1.525 ;
        RECT 428.235 1.195 428.565 1.525 ;
        RECT 426.875 1.195 427.205 1.525 ;
        RECT 425.515 1.195 425.845 1.525 ;
        RECT 424.155 1.195 424.485 1.525 ;
        RECT 422.795 1.195 423.125 1.525 ;
        RECT 421.435 1.195 421.765 1.525 ;
        RECT 420.075 1.195 420.405 1.525 ;
        RECT 418.715 1.195 419.045 1.525 ;
        RECT 417.355 1.195 417.685 1.525 ;
        RECT 415.995 1.195 416.325 1.525 ;
        RECT 414.635 1.195 414.965 1.525 ;
        RECT 413.275 1.195 413.605 1.525 ;
        RECT 411.915 1.195 412.245 1.525 ;
        RECT 410.555 1.195 410.885 1.525 ;
        RECT 409.195 1.195 409.525 1.525 ;
        RECT 407.835 1.195 408.165 1.525 ;
        RECT 406.475 1.195 406.805 1.525 ;
        RECT 405.115 1.195 405.445 1.525 ;
        RECT 403.755 1.195 404.085 1.525 ;
        RECT 402.395 1.195 402.725 1.525 ;
        RECT 401.035 1.195 401.365 1.525 ;
        RECT 399.675 1.195 400.005 1.525 ;
        RECT 398.315 1.195 398.645 1.525 ;
        RECT 396.955 1.195 397.285 1.525 ;
        RECT 395.595 1.195 395.925 1.525 ;
        RECT 394.235 1.195 394.565 1.525 ;
        RECT 392.875 1.195 393.205 1.525 ;
        RECT 391.515 1.195 391.845 1.525 ;
        RECT 390.155 1.195 390.485 1.525 ;
        RECT 388.795 1.195 389.125 1.525 ;
        RECT 387.435 1.195 387.765 1.525 ;
        RECT 386.075 1.195 386.405 1.525 ;
        RECT 384.715 1.195 385.045 1.525 ;
        RECT 383.355 1.195 383.685 1.525 ;
        RECT 381.995 1.195 382.325 1.525 ;
        RECT 380.635 1.195 380.965 1.525 ;
        RECT 379.275 1.195 379.605 1.525 ;
        RECT 377.915 1.195 378.245 1.525 ;
        RECT 376.555 1.195 376.885 1.525 ;
        RECT 375.195 1.195 375.525 1.525 ;
        RECT 373.835 1.195 374.165 1.525 ;
        RECT 372.475 1.195 372.805 1.525 ;
        RECT 371.115 1.195 371.445 1.525 ;
        RECT 369.755 1.195 370.085 1.525 ;
        RECT 368.395 1.195 368.725 1.525 ;
        RECT 367.035 1.195 367.365 1.525 ;
        RECT 365.675 1.195 366.005 1.525 ;
        RECT 364.315 1.195 364.645 1.525 ;
        RECT 362.955 1.195 363.285 1.525 ;
        RECT 361.595 1.195 361.925 1.525 ;
        RECT 360.235 1.195 360.565 1.525 ;
        RECT 358.875 1.195 359.205 1.525 ;
        RECT 357.515 1.195 357.845 1.525 ;
        RECT 356.155 1.195 356.485 1.525 ;
        RECT 354.795 1.195 355.125 1.525 ;
        RECT 353.435 1.195 353.765 1.525 ;
        RECT 352.075 1.195 352.405 1.525 ;
        RECT 350.715 1.195 351.045 1.525 ;
        RECT 349.355 1.195 349.685 1.525 ;
        RECT 347.995 1.195 348.325 1.525 ;
        RECT 346.635 1.195 346.965 1.525 ;
        RECT 345.275 1.195 345.605 1.525 ;
        RECT 343.915 1.195 344.245 1.525 ;
        RECT 342.555 1.195 342.885 1.525 ;
        RECT 341.195 1.195 341.525 1.525 ;
        RECT 339.835 1.195 340.165 1.525 ;
        RECT 338.475 1.195 338.805 1.525 ;
        RECT 337.115 1.195 337.445 1.525 ;
        RECT 335.755 1.195 336.085 1.525 ;
        RECT 334.395 1.195 334.725 1.525 ;
        RECT 333.035 1.195 333.365 1.525 ;
        RECT 331.675 1.195 332.005 1.525 ;
        RECT 330.315 1.195 330.645 1.525 ;
        RECT 328.955 1.195 329.285 1.525 ;
        RECT 327.595 1.195 327.925 1.525 ;
        RECT 326.235 1.195 326.565 1.525 ;
        RECT 324.875 1.195 325.205 1.525 ;
        RECT 323.515 1.195 323.845 1.525 ;
        RECT 322.155 1.195 322.485 1.525 ;
        RECT 320.795 1.195 321.125 1.525 ;
        RECT 319.435 1.195 319.765 1.525 ;
        RECT 318.075 1.195 318.405 1.525 ;
        RECT 316.715 1.195 317.045 1.525 ;
        RECT 315.355 1.195 315.685 1.525 ;
        RECT 313.995 1.195 314.325 1.525 ;
        RECT 312.635 1.195 312.965 1.525 ;
        RECT 311.275 1.195 311.605 1.525 ;
        RECT 309.915 1.195 310.245 1.525 ;
        RECT 308.555 1.195 308.885 1.525 ;
        RECT 307.195 1.195 307.525 1.525 ;
        RECT 305.835 1.195 306.165 1.525 ;
        RECT 304.475 1.195 304.805 1.525 ;
        RECT 303.115 1.195 303.445 1.525 ;
        RECT 301.755 1.195 302.085 1.525 ;
        RECT 300.395 1.195 300.725 1.525 ;
        RECT 299.035 1.195 299.365 1.525 ;
        RECT 297.675 1.195 298.005 1.525 ;
        RECT 296.315 1.195 296.645 1.525 ;
        RECT 294.955 1.195 295.285 1.525 ;
        RECT 293.595 1.195 293.925 1.525 ;
        RECT 292.235 1.195 292.565 1.525 ;
        RECT 290.875 1.195 291.205 1.525 ;
        RECT 289.515 1.195 289.845 1.525 ;
        RECT 288.155 1.195 288.485 1.525 ;
        RECT 286.795 1.195 287.125 1.525 ;
        RECT 285.435 1.195 285.765 1.525 ;
        RECT 284.075 1.195 284.405 1.525 ;
        RECT 282.715 1.195 283.045 1.525 ;
        RECT 281.355 1.195 281.685 1.525 ;
        RECT 279.995 1.195 280.325 1.525 ;
        RECT 278.635 1.195 278.965 1.525 ;
        RECT 277.275 1.195 277.605 1.525 ;
        RECT 275.915 1.195 276.245 1.525 ;
        RECT 274.555 1.195 274.885 1.525 ;
        RECT 273.195 1.195 273.525 1.525 ;
        RECT 271.835 1.195 272.165 1.525 ;
        RECT 270.475 1.195 270.805 1.525 ;
        RECT 269.115 1.195 269.445 1.525 ;
        RECT 267.755 1.195 268.085 1.525 ;
        RECT 266.395 1.195 266.725 1.525 ;
        RECT 265.035 1.195 265.365 1.525 ;
        RECT 263.675 1.195 264.005 1.525 ;
        RECT 262.315 1.195 262.645 1.525 ;
        RECT 260.955 1.195 261.285 1.525 ;
        RECT 259.595 1.195 259.925 1.525 ;
        RECT 258.235 1.195 258.565 1.525 ;
        RECT 256.875 1.195 257.205 1.525 ;
        RECT 255.515 1.195 255.845 1.525 ;
        RECT 254.155 1.195 254.485 1.525 ;
        RECT 252.795 1.195 253.125 1.525 ;
        RECT 251.435 1.195 251.765 1.525 ;
        RECT 250.075 1.195 250.405 1.525 ;
        RECT 248.715 1.195 249.045 1.525 ;
        RECT 247.355 1.195 247.685 1.525 ;
        RECT 245.995 1.195 246.325 1.525 ;
        RECT 244.635 1.195 244.965 1.525 ;
        RECT 243.275 1.195 243.605 1.525 ;
        RECT 241.915 1.195 242.245 1.525 ;
        RECT 240.555 1.195 240.885 1.525 ;
        RECT 239.195 1.195 239.525 1.525 ;
        RECT 237.835 1.195 238.165 1.525 ;
        RECT 236.475 1.195 236.805 1.525 ;
        RECT 235.115 1.195 235.445 1.525 ;
        RECT 233.755 1.195 234.085 1.525 ;
        RECT 232.395 1.195 232.725 1.525 ;
        RECT 231.035 1.195 231.365 1.525 ;
        RECT 229.675 1.195 230.005 1.525 ;
        RECT 228.315 1.195 228.645 1.525 ;
        RECT 226.955 1.195 227.285 1.525 ;
        RECT 225.595 1.195 225.925 1.525 ;
        RECT 224.235 1.195 224.565 1.525 ;
        RECT 222.875 1.195 223.205 1.525 ;
        RECT 221.515 1.195 221.845 1.525 ;
        RECT 220.155 1.195 220.485 1.525 ;
        RECT 218.795 1.195 219.125 1.525 ;
        RECT 217.435 1.195 217.765 1.525 ;
        RECT 216.075 1.195 216.405 1.525 ;
        RECT 214.715 1.195 215.045 1.525 ;
        RECT 213.355 1.195 213.685 1.525 ;
        RECT 211.995 1.195 212.325 1.525 ;
        RECT 210.635 1.195 210.965 1.525 ;
        RECT 209.275 1.195 209.605 1.525 ;
        RECT 207.915 1.195 208.245 1.525 ;
        RECT 206.555 1.195 206.885 1.525 ;
        RECT 205.195 1.195 205.525 1.525 ;
        RECT 203.835 1.195 204.165 1.525 ;
        RECT 202.475 1.195 202.805 1.525 ;
        RECT 201.115 1.195 201.445 1.525 ;
        RECT 199.755 1.195 200.085 1.525 ;
        RECT 198.395 1.195 198.725 1.525 ;
        RECT 197.035 1.195 197.365 1.525 ;
        RECT 195.675 1.195 196.005 1.525 ;
        RECT 194.315 1.195 194.645 1.525 ;
        RECT 192.955 1.195 193.285 1.525 ;
        RECT 191.595 1.195 191.925 1.525 ;
        RECT 190.235 1.195 190.565 1.525 ;
        RECT 188.875 1.195 189.205 1.525 ;
        RECT 187.515 1.195 187.845 1.525 ;
        RECT 186.155 1.195 186.485 1.525 ;
        RECT 184.795 1.195 185.125 1.525 ;
        RECT 183.435 1.195 183.765 1.525 ;
        RECT 182.075 1.195 182.405 1.525 ;
        RECT 180.715 1.195 181.045 1.525 ;
        RECT 179.355 1.195 179.685 1.525 ;
        RECT 177.995 1.195 178.325 1.525 ;
        RECT 176.635 1.195 176.965 1.525 ;
        RECT 175.275 1.195 175.605 1.525 ;
        RECT 173.915 1.195 174.245 1.525 ;
        RECT 172.555 1.195 172.885 1.525 ;
        RECT 171.195 1.195 171.525 1.525 ;
        RECT 169.835 1.195 170.165 1.525 ;
        RECT 168.475 1.195 168.805 1.525 ;
        RECT 167.115 1.195 167.445 1.525 ;
        RECT 165.755 1.195 166.085 1.525 ;
        RECT 164.395 1.195 164.725 1.525 ;
        RECT 163.035 1.195 163.365 1.525 ;
        RECT 161.675 1.195 162.005 1.525 ;
        RECT 160.315 1.195 160.645 1.525 ;
        RECT 158.955 1.195 159.285 1.525 ;
        RECT 157.595 1.195 157.925 1.525 ;
        RECT 156.235 1.195 156.565 1.525 ;
        RECT 154.875 1.195 155.205 1.525 ;
        RECT 153.515 1.195 153.845 1.525 ;
        RECT 152.155 1.195 152.485 1.525 ;
        RECT 150.795 1.195 151.125 1.525 ;
        RECT 149.435 1.195 149.765 1.525 ;
        RECT 148.075 1.195 148.405 1.525 ;
        RECT 146.715 1.195 147.045 1.525 ;
        RECT 145.355 1.195 145.685 1.525 ;
        RECT 143.995 1.195 144.325 1.525 ;
        RECT 142.635 1.195 142.965 1.525 ;
        RECT 141.275 1.195 141.605 1.525 ;
        RECT 139.915 1.195 140.245 1.525 ;
        RECT 138.555 1.195 138.885 1.525 ;
        RECT 137.195 1.195 137.525 1.525 ;
        RECT 135.835 1.195 136.165 1.525 ;
        RECT 134.475 1.195 134.805 1.525 ;
        RECT 133.115 1.195 133.445 1.525 ;
        RECT 131.755 1.195 132.085 1.525 ;
        RECT 130.395 1.195 130.725 1.525 ;
        RECT 129.035 1.195 129.365 1.525 ;
        RECT 127.675 1.195 128.005 1.525 ;
        RECT 126.315 1.195 126.645 1.525 ;
        RECT 124.955 1.195 125.285 1.525 ;
        RECT 123.595 1.195 123.925 1.525 ;
        RECT 122.235 1.195 122.565 1.525 ;
        RECT 120.875 1.195 121.205 1.525 ;
        RECT 119.515 1.195 119.845 1.525 ;
        RECT 118.155 1.195 118.485 1.525 ;
        RECT 116.795 1.195 117.125 1.525 ;
        RECT 115.435 1.195 115.765 1.525 ;
        RECT 114.075 1.195 114.405 1.525 ;
        RECT 112.715 1.195 113.045 1.525 ;
        RECT 111.355 1.195 111.685 1.525 ;
        RECT 109.995 1.195 110.325 1.525 ;
        RECT 108.635 1.195 108.965 1.525 ;
        RECT 107.275 1.195 107.605 1.525 ;
        RECT 105.915 1.195 106.245 1.525 ;
        RECT 104.555 1.195 104.885 1.525 ;
        RECT 103.195 1.195 103.525 1.525 ;
        RECT 101.835 1.195 102.165 1.525 ;
        RECT 100.475 1.195 100.805 1.525 ;
        RECT 99.115 1.195 99.445 1.525 ;
        RECT 97.755 1.195 98.085 1.525 ;
        RECT 96.395 1.195 96.725 1.525 ;
        RECT 95.035 1.195 95.365 1.525 ;
        RECT 93.675 1.195 94.005 1.525 ;
        RECT 92.315 1.195 92.645 1.525 ;
        RECT 90.955 1.195 91.285 1.525 ;
        RECT 89.595 1.195 89.925 1.525 ;
        RECT 88.235 1.195 88.565 1.525 ;
        RECT 86.875 1.195 87.205 1.525 ;
        RECT 85.515 1.195 85.845 1.525 ;
        RECT 84.155 1.195 84.485 1.525 ;
        RECT 82.795 1.195 83.125 1.525 ;
        RECT 81.435 1.195 81.765 1.525 ;
        RECT 80.075 1.195 80.405 1.525 ;
        RECT 78.715 1.195 79.045 1.525 ;
        RECT 77.355 1.195 77.685 1.525 ;
        RECT 75.995 1.195 76.325 1.525 ;
        RECT 74.635 1.195 74.965 1.525 ;
        RECT 73.275 1.195 73.605 1.525 ;
        RECT 71.915 1.195 72.245 1.525 ;
        RECT 70.555 1.195 70.885 1.525 ;
        RECT 69.195 1.195 69.525 1.525 ;
        RECT 67.835 1.195 68.165 1.525 ;
        RECT 66.475 1.195 66.805 1.525 ;
        RECT 65.115 1.195 65.445 1.525 ;
        RECT 63.755 1.195 64.085 1.525 ;
        RECT 62.395 1.195 62.725 1.525 ;
        RECT 61.035 1.195 61.365 1.525 ;
        RECT 59.675 1.195 60.005 1.525 ;
        RECT 58.315 1.195 58.645 1.525 ;
        RECT 56.955 1.195 57.285 1.525 ;
        RECT 55.595 1.195 55.925 1.525 ;
        RECT 54.235 1.195 54.565 1.525 ;
        RECT 52.875 1.195 53.205 1.525 ;
        RECT 51.515 1.195 51.845 1.525 ;
        RECT 50.155 1.195 50.485 1.525 ;
        RECT 48.795 1.195 49.125 1.525 ;
        RECT 47.435 1.195 47.765 1.525 ;
        RECT 46.075 1.195 46.405 1.525 ;
        RECT 44.715 1.195 45.045 1.525 ;
        RECT 43.355 1.195 43.685 1.525 ;
        RECT 41.995 1.195 42.325 1.525 ;
        RECT 40.635 1.195 40.965 1.525 ;
        RECT 39.275 1.195 39.605 1.525 ;
        RECT 37.915 1.195 38.245 1.525 ;
        RECT 36.555 1.195 36.885 1.525 ;
        RECT 35.195 1.195 35.525 1.525 ;
        RECT 33.835 1.195 34.165 1.525 ;
        RECT 32.475 1.195 32.805 1.525 ;
        RECT 31.115 1.195 31.445 1.525 ;
        RECT 29.755 1.195 30.085 1.525 ;
        RECT 28.395 1.195 28.725 1.525 ;
        RECT 27.035 1.195 27.365 1.525 ;
        RECT 25.675 1.195 26.005 1.525 ;
        RECT 24.315 1.195 24.645 1.525 ;
        RECT 22.955 1.195 23.285 1.525 ;
        RECT 21.595 1.195 21.925 1.525 ;
        RECT 20.235 1.195 20.565 1.525 ;
        RECT 18.875 1.195 19.205 1.525 ;
        RECT 17.515 1.195 17.845 1.525 ;
        RECT 16.155 1.195 16.485 1.525 ;
        RECT 14.795 1.195 15.125 1.525 ;
        RECT 13.435 1.195 13.765 1.525 ;
        RECT 12.075 1.195 12.405 1.525 ;
        RECT 10.715 1.195 11.045 1.525 ;
        RECT 9.355 1.195 9.685 1.525 ;
        RECT 7.995 1.195 8.325 1.525 ;
        RECT 6.635 1.195 6.965 1.525 ;
        RECT 5.275 1.195 5.605 1.525 ;
        RECT 3.915 1.195 4.245 1.525 ;
        RECT 2.555 1.195 2.885 1.525 ;
        RECT 1.195 1.195 1.525 1.525 ;
        RECT -0.165 1.195 0.165 1.525 ;
        RECT -1.525 1.195 -1.195 1.525 ;
        RECT 954.555 1.195 954.885 1.525 ;
        RECT 678.475 1.2 954.885 1.52 ;
        RECT 953.195 1.195 953.525 1.525 ;
        RECT 951.835 1.195 952.165 1.525 ;
        RECT 950.475 1.195 950.805 1.525 ;
        RECT 949.115 1.195 949.445 1.525 ;
        RECT 947.755 1.195 948.085 1.525 ;
        RECT 946.395 1.195 946.725 1.525 ;
        RECT 945.035 1.195 945.365 1.525 ;
        RECT 943.675 1.195 944.005 1.525 ;
        RECT 942.315 1.195 942.645 1.525 ;
        RECT 940.955 1.195 941.285 1.525 ;
        RECT 939.595 1.195 939.925 1.525 ;
        RECT 938.235 1.195 938.565 1.525 ;
        RECT 936.875 1.195 937.205 1.525 ;
        RECT 935.515 1.195 935.845 1.525 ;
        RECT 934.155 1.195 934.485 1.525 ;
        RECT 932.795 1.195 933.125 1.525 ;
        RECT 931.435 1.195 931.765 1.525 ;
        RECT 930.075 1.195 930.405 1.525 ;
        RECT 928.715 1.195 929.045 1.525 ;
        RECT 927.355 1.195 927.685 1.525 ;
        RECT 925.995 1.195 926.325 1.525 ;
        RECT 924.635 1.195 924.965 1.525 ;
        RECT 923.275 1.195 923.605 1.525 ;
        RECT 921.915 1.195 922.245 1.525 ;
        RECT 920.555 1.195 920.885 1.525 ;
        RECT 919.195 1.195 919.525 1.525 ;
        RECT 917.835 1.195 918.165 1.525 ;
        RECT 916.475 1.195 916.805 1.525 ;
        RECT 915.115 1.195 915.445 1.525 ;
        RECT 913.755 1.195 914.085 1.525 ;
        RECT 912.395 1.195 912.725 1.525 ;
        RECT 911.035 1.195 911.365 1.525 ;
        RECT 909.675 1.195 910.005 1.525 ;
        RECT 908.315 1.195 908.645 1.525 ;
        RECT 906.955 1.195 907.285 1.525 ;
        RECT 905.595 1.195 905.925 1.525 ;
        RECT 904.235 1.195 904.565 1.525 ;
        RECT 902.875 1.195 903.205 1.525 ;
        RECT 901.515 1.195 901.845 1.525 ;
        RECT 900.155 1.195 900.485 1.525 ;
        RECT 898.795 1.195 899.125 1.525 ;
        RECT 897.435 1.195 897.765 1.525 ;
        RECT 896.075 1.195 896.405 1.525 ;
        RECT 894.715 1.195 895.045 1.525 ;
        RECT 893.355 1.195 893.685 1.525 ;
        RECT 891.995 1.195 892.325 1.525 ;
        RECT 890.635 1.195 890.965 1.525 ;
        RECT 889.275 1.195 889.605 1.525 ;
        RECT 887.915 1.195 888.245 1.525 ;
        RECT 886.555 1.195 886.885 1.525 ;
        RECT 885.195 1.195 885.525 1.525 ;
        RECT 883.835 1.195 884.165 1.525 ;
        RECT 882.475 1.195 882.805 1.525 ;
        RECT 881.115 1.195 881.445 1.525 ;
        RECT 879.755 1.195 880.085 1.525 ;
        RECT 878.395 1.195 878.725 1.525 ;
        RECT 877.035 1.195 877.365 1.525 ;
        RECT 875.675 1.195 876.005 1.525 ;
        RECT 874.315 1.195 874.645 1.525 ;
        RECT 872.955 1.195 873.285 1.525 ;
        RECT 871.595 1.195 871.925 1.525 ;
        RECT 870.235 1.195 870.565 1.525 ;
        RECT 868.875 1.195 869.205 1.525 ;
        RECT 867.515 1.195 867.845 1.525 ;
        RECT 866.155 1.195 866.485 1.525 ;
        RECT 864.795 1.195 865.125 1.525 ;
        RECT 863.435 1.195 863.765 1.525 ;
        RECT 862.075 1.195 862.405 1.525 ;
        RECT 860.715 1.195 861.045 1.525 ;
        RECT 859.355 1.195 859.685 1.525 ;
        RECT 857.995 1.195 858.325 1.525 ;
        RECT 856.635 1.195 856.965 1.525 ;
        RECT 855.275 1.195 855.605 1.525 ;
        RECT 853.915 1.195 854.245 1.525 ;
        RECT 852.555 1.195 852.885 1.525 ;
        RECT 851.195 1.195 851.525 1.525 ;
        RECT 849.835 1.195 850.165 1.525 ;
        RECT 848.475 1.195 848.805 1.525 ;
        RECT 847.115 1.195 847.445 1.525 ;
        RECT 845.755 1.195 846.085 1.525 ;
        RECT 844.395 1.195 844.725 1.525 ;
        RECT 843.035 1.195 843.365 1.525 ;
        RECT 841.675 1.195 842.005 1.525 ;
        RECT 840.315 1.195 840.645 1.525 ;
        RECT 838.955 1.195 839.285 1.525 ;
        RECT 837.595 1.195 837.925 1.525 ;
        RECT 836.235 1.195 836.565 1.525 ;
        RECT 834.875 1.195 835.205 1.525 ;
        RECT 833.515 1.195 833.845 1.525 ;
        RECT 832.155 1.195 832.485 1.525 ;
        RECT 830.795 1.195 831.125 1.525 ;
        RECT 829.435 1.195 829.765 1.525 ;
        RECT 828.075 1.195 828.405 1.525 ;
        RECT 826.715 1.195 827.045 1.525 ;
        RECT 825.355 1.195 825.685 1.525 ;
        RECT 823.995 1.195 824.325 1.525 ;
        RECT 822.635 1.195 822.965 1.525 ;
        RECT 821.275 1.195 821.605 1.525 ;
        RECT 819.915 1.195 820.245 1.525 ;
        RECT 818.555 1.195 818.885 1.525 ;
        RECT 817.195 1.195 817.525 1.525 ;
        RECT 815.835 1.195 816.165 1.525 ;
        RECT 814.475 1.195 814.805 1.525 ;
        RECT 813.115 1.195 813.445 1.525 ;
        RECT 811.755 1.195 812.085 1.525 ;
        RECT 810.395 1.195 810.725 1.525 ;
        RECT 809.035 1.195 809.365 1.525 ;
        RECT 807.675 1.195 808.005 1.525 ;
        RECT 806.315 1.195 806.645 1.525 ;
        RECT 804.955 1.195 805.285 1.525 ;
        RECT 803.595 1.195 803.925 1.525 ;
        RECT 802.235 1.195 802.565 1.525 ;
        RECT 800.875 1.195 801.205 1.525 ;
        RECT 799.515 1.195 799.845 1.525 ;
        RECT 798.155 1.195 798.485 1.525 ;
        RECT 796.795 1.195 797.125 1.525 ;
        RECT 795.435 1.195 795.765 1.525 ;
        RECT 794.075 1.195 794.405 1.525 ;
        RECT 792.715 1.195 793.045 1.525 ;
        RECT 791.355 1.195 791.685 1.525 ;
        RECT 789.995 1.195 790.325 1.525 ;
        RECT 788.635 1.195 788.965 1.525 ;
        RECT 787.275 1.195 787.605 1.525 ;
        RECT 785.915 1.195 786.245 1.525 ;
        RECT 784.555 1.195 784.885 1.525 ;
        RECT 783.195 1.195 783.525 1.525 ;
        RECT 781.835 1.195 782.165 1.525 ;
        RECT 780.475 1.195 780.805 1.525 ;
        RECT 779.115 1.195 779.445 1.525 ;
        RECT 777.755 1.195 778.085 1.525 ;
        RECT 776.395 1.195 776.725 1.525 ;
        RECT 775.035 1.195 775.365 1.525 ;
        RECT 773.675 1.195 774.005 1.525 ;
        RECT 772.315 1.195 772.645 1.525 ;
        RECT 770.955 1.195 771.285 1.525 ;
        RECT 769.595 1.195 769.925 1.525 ;
        RECT 768.235 1.195 768.565 1.525 ;
        RECT 766.875 1.195 767.205 1.525 ;
        RECT 765.515 1.195 765.845 1.525 ;
        RECT 764.155 1.195 764.485 1.525 ;
        RECT 762.795 1.195 763.125 1.525 ;
        RECT 761.435 1.195 761.765 1.525 ;
        RECT 760.075 1.195 760.405 1.525 ;
        RECT 758.715 1.195 759.045 1.525 ;
        RECT 757.355 1.195 757.685 1.525 ;
        RECT 755.995 1.195 756.325 1.525 ;
        RECT 754.635 1.195 754.965 1.525 ;
        RECT 753.275 1.195 753.605 1.525 ;
        RECT 751.915 1.195 752.245 1.525 ;
        RECT 750.555 1.195 750.885 1.525 ;
        RECT 749.195 1.195 749.525 1.525 ;
        RECT 747.835 1.195 748.165 1.525 ;
        RECT 746.475 1.195 746.805 1.525 ;
        RECT 745.115 1.195 745.445 1.525 ;
        RECT 743.755 1.195 744.085 1.525 ;
        RECT 742.395 1.195 742.725 1.525 ;
        RECT 741.035 1.195 741.365 1.525 ;
        RECT 739.675 1.195 740.005 1.525 ;
        RECT 738.315 1.195 738.645 1.525 ;
        RECT 736.955 1.195 737.285 1.525 ;
        RECT 735.595 1.195 735.925 1.525 ;
        RECT 734.235 1.195 734.565 1.525 ;
        RECT 732.875 1.195 733.205 1.525 ;
        RECT 731.515 1.195 731.845 1.525 ;
        RECT 730.155 1.195 730.485 1.525 ;
        RECT 728.795 1.195 729.125 1.525 ;
        RECT 727.435 1.195 727.765 1.525 ;
        RECT 726.075 1.195 726.405 1.525 ;
        RECT 724.715 1.195 725.045 1.525 ;
        RECT 723.355 1.195 723.685 1.525 ;
        RECT 721.995 1.195 722.325 1.525 ;
        RECT 720.635 1.195 720.965 1.525 ;
        RECT 719.275 1.195 719.605 1.525 ;
        RECT 717.915 1.195 718.245 1.525 ;
        RECT 716.555 1.195 716.885 1.525 ;
        RECT 715.195 1.195 715.525 1.525 ;
        RECT 713.835 1.195 714.165 1.525 ;
        RECT 712.475 1.195 712.805 1.525 ;
        RECT 711.115 1.195 711.445 1.525 ;
        RECT 709.755 1.195 710.085 1.525 ;
        RECT 708.395 1.195 708.725 1.525 ;
        RECT 707.035 1.195 707.365 1.525 ;
        RECT 705.675 1.195 706.005 1.525 ;
        RECT 704.315 1.195 704.645 1.525 ;
        RECT 702.955 1.195 703.285 1.525 ;
        RECT 701.595 1.195 701.925 1.525 ;
        RECT 700.235 1.195 700.565 1.525 ;
        RECT 698.875 1.195 699.205 1.525 ;
        RECT 697.515 1.195 697.845 1.525 ;
        RECT 696.155 1.195 696.485 1.525 ;
        RECT 694.795 1.195 695.125 1.525 ;
        RECT 693.435 1.195 693.765 1.525 ;
        RECT 692.075 1.195 692.405 1.525 ;
        RECT 690.715 1.195 691.045 1.525 ;
        RECT 689.355 1.195 689.685 1.525 ;
        RECT 687.995 1.195 688.325 1.525 ;
        RECT 686.635 1.195 686.965 1.525 ;
        RECT 685.275 1.195 685.605 1.525 ;
        RECT 683.915 1.195 684.245 1.525 ;
        RECT 682.555 1.195 682.885 1.525 ;
        RECT 681.195 1.195 681.525 1.525 ;
        RECT 679.835 1.195 680.165 1.525 ;
        RECT 678.475 1.195 678.805 1.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 659.435 -0.165 659.765 0.165 ;
        RECT 658.075 -0.165 658.405 0.165 ;
        RECT 656.715 -0.165 657.045 0.165 ;
        RECT 655.355 -0.165 655.685 0.165 ;
        RECT 653.995 -0.165 654.325 0.165 ;
        RECT 652.635 -0.165 652.965 0.165 ;
        RECT 651.275 -0.165 651.605 0.165 ;
        RECT 649.915 -0.165 650.245 0.165 ;
        RECT 648.555 -0.165 648.885 0.165 ;
        RECT 647.195 -0.165 647.525 0.165 ;
        RECT 645.835 -0.165 646.165 0.165 ;
        RECT 644.475 -0.165 644.805 0.165 ;
        RECT 643.115 -0.165 643.445 0.165 ;
        RECT 641.755 -0.165 642.085 0.165 ;
        RECT 640.395 -0.165 640.725 0.165 ;
        RECT 639.035 -0.165 639.365 0.165 ;
        RECT 637.675 -0.165 638.005 0.165 ;
        RECT 636.315 -0.165 636.645 0.165 ;
        RECT 634.955 -0.165 635.285 0.165 ;
        RECT 633.595 -0.165 633.925 0.165 ;
        RECT 632.235 -0.165 632.565 0.165 ;
        RECT 630.875 -0.165 631.205 0.165 ;
        RECT 629.515 -0.165 629.845 0.165 ;
        RECT 628.155 -0.165 628.485 0.165 ;
        RECT 626.795 -0.165 627.125 0.165 ;
        RECT 625.435 -0.165 625.765 0.165 ;
        RECT 624.075 -0.165 624.405 0.165 ;
        RECT 622.715 -0.165 623.045 0.165 ;
        RECT 621.355 -0.165 621.685 0.165 ;
        RECT 619.995 -0.165 620.325 0.165 ;
        RECT 618.635 -0.165 618.965 0.165 ;
        RECT 617.275 -0.165 617.605 0.165 ;
        RECT 615.915 -0.165 616.245 0.165 ;
        RECT 614.555 -0.165 614.885 0.165 ;
        RECT 613.195 -0.165 613.525 0.165 ;
        RECT 611.835 -0.165 612.165 0.165 ;
        RECT 610.475 -0.165 610.805 0.165 ;
        RECT 609.115 -0.165 609.445 0.165 ;
        RECT 607.755 -0.165 608.085 0.165 ;
        RECT 606.395 -0.165 606.725 0.165 ;
        RECT 605.035 -0.165 605.365 0.165 ;
        RECT 603.675 -0.165 604.005 0.165 ;
        RECT 602.315 -0.165 602.645 0.165 ;
        RECT 600.955 -0.165 601.285 0.165 ;
        RECT 599.595 -0.165 599.925 0.165 ;
        RECT 598.235 -0.165 598.565 0.165 ;
        RECT 596.875 -0.165 597.205 0.165 ;
        RECT 595.515 -0.165 595.845 0.165 ;
        RECT 594.155 -0.165 594.485 0.165 ;
        RECT 592.795 -0.165 593.125 0.165 ;
        RECT 591.435 -0.165 591.765 0.165 ;
        RECT 590.075 -0.165 590.405 0.165 ;
        RECT 588.715 -0.165 589.045 0.165 ;
        RECT 587.355 -0.165 587.685 0.165 ;
        RECT 585.995 -0.165 586.325 0.165 ;
        RECT 584.635 -0.165 584.965 0.165 ;
        RECT 583.275 -0.165 583.605 0.165 ;
        RECT 581.915 -0.165 582.245 0.165 ;
        RECT 580.555 -0.165 580.885 0.165 ;
        RECT 579.195 -0.165 579.525 0.165 ;
        RECT 577.835 -0.165 578.165 0.165 ;
        RECT 576.475 -0.165 576.805 0.165 ;
        RECT 575.115 -0.165 575.445 0.165 ;
        RECT 573.755 -0.165 574.085 0.165 ;
        RECT 572.395 -0.165 572.725 0.165 ;
        RECT 571.035 -0.165 571.365 0.165 ;
        RECT 569.675 -0.165 570.005 0.165 ;
        RECT 568.315 -0.165 568.645 0.165 ;
        RECT 566.955 -0.165 567.285 0.165 ;
        RECT 565.595 -0.165 565.925 0.165 ;
        RECT 564.235 -0.165 564.565 0.165 ;
        RECT 562.875 -0.165 563.205 0.165 ;
        RECT 561.515 -0.165 561.845 0.165 ;
        RECT 560.155 -0.165 560.485 0.165 ;
        RECT 558.795 -0.165 559.125 0.165 ;
        RECT 557.435 -0.165 557.765 0.165 ;
        RECT 556.075 -0.165 556.405 0.165 ;
        RECT 554.715 -0.165 555.045 0.165 ;
        RECT 553.355 -0.165 553.685 0.165 ;
        RECT 551.995 -0.165 552.325 0.165 ;
        RECT 550.635 -0.165 550.965 0.165 ;
        RECT 549.275 -0.165 549.605 0.165 ;
        RECT 547.915 -0.165 548.245 0.165 ;
        RECT 546.555 -0.165 546.885 0.165 ;
        RECT 545.195 -0.165 545.525 0.165 ;
        RECT 543.835 -0.165 544.165 0.165 ;
        RECT 542.475 -0.165 542.805 0.165 ;
        RECT 541.115 -0.165 541.445 0.165 ;
        RECT 539.755 -0.165 540.085 0.165 ;
        RECT 538.395 -0.165 538.725 0.165 ;
        RECT 537.035 -0.165 537.365 0.165 ;
        RECT 535.675 -0.165 536.005 0.165 ;
        RECT 534.315 -0.165 534.645 0.165 ;
        RECT 532.955 -0.165 533.285 0.165 ;
        RECT 531.595 -0.165 531.925 0.165 ;
        RECT 530.235 -0.165 530.565 0.165 ;
        RECT 528.875 -0.165 529.205 0.165 ;
        RECT 527.515 -0.165 527.845 0.165 ;
        RECT 526.155 -0.165 526.485 0.165 ;
        RECT 524.795 -0.165 525.125 0.165 ;
        RECT 523.435 -0.165 523.765 0.165 ;
        RECT 522.075 -0.165 522.405 0.165 ;
        RECT 520.715 -0.165 521.045 0.165 ;
        RECT 519.355 -0.165 519.685 0.165 ;
        RECT 517.995 -0.165 518.325 0.165 ;
        RECT 516.635 -0.165 516.965 0.165 ;
        RECT 515.275 -0.165 515.605 0.165 ;
        RECT 513.915 -0.165 514.245 0.165 ;
        RECT 512.555 -0.165 512.885 0.165 ;
        RECT 511.195 -0.165 511.525 0.165 ;
        RECT 509.835 -0.165 510.165 0.165 ;
        RECT 508.475 -0.165 508.805 0.165 ;
        RECT 507.115 -0.165 507.445 0.165 ;
        RECT 505.755 -0.165 506.085 0.165 ;
        RECT 504.395 -0.165 504.725 0.165 ;
        RECT 503.035 -0.165 503.365 0.165 ;
        RECT 501.675 -0.165 502.005 0.165 ;
        RECT 500.315 -0.165 500.645 0.165 ;
        RECT 498.955 -0.165 499.285 0.165 ;
        RECT 497.595 -0.165 497.925 0.165 ;
        RECT 496.235 -0.165 496.565 0.165 ;
        RECT 494.875 -0.165 495.205 0.165 ;
        RECT 493.515 -0.165 493.845 0.165 ;
        RECT 492.155 -0.165 492.485 0.165 ;
        RECT 490.795 -0.165 491.125 0.165 ;
        RECT 489.435 -0.165 489.765 0.165 ;
        RECT 488.075 -0.165 488.405 0.165 ;
        RECT 486.715 -0.165 487.045 0.165 ;
        RECT 485.355 -0.165 485.685 0.165 ;
        RECT 483.995 -0.165 484.325 0.165 ;
        RECT 482.635 -0.165 482.965 0.165 ;
        RECT 481.275 -0.165 481.605 0.165 ;
        RECT 479.915 -0.165 480.245 0.165 ;
        RECT 478.555 -0.165 478.885 0.165 ;
        RECT 477.195 -0.165 477.525 0.165 ;
        RECT 475.835 -0.165 476.165 0.165 ;
        RECT 474.475 -0.165 474.805 0.165 ;
        RECT 473.115 -0.165 473.445 0.165 ;
        RECT 471.755 -0.165 472.085 0.165 ;
        RECT 470.395 -0.165 470.725 0.165 ;
        RECT 469.035 -0.165 469.365 0.165 ;
        RECT 467.675 -0.165 468.005 0.165 ;
        RECT 466.315 -0.165 466.645 0.165 ;
        RECT 464.955 -0.165 465.285 0.165 ;
        RECT 463.595 -0.165 463.925 0.165 ;
        RECT 462.235 -0.165 462.565 0.165 ;
        RECT 460.875 -0.165 461.205 0.165 ;
        RECT 459.515 -0.165 459.845 0.165 ;
        RECT 458.155 -0.165 458.485 0.165 ;
        RECT 456.795 -0.165 457.125 0.165 ;
        RECT 455.435 -0.165 455.765 0.165 ;
        RECT 454.075 -0.165 454.405 0.165 ;
        RECT 452.715 -0.165 453.045 0.165 ;
        RECT 451.355 -0.165 451.685 0.165 ;
        RECT 449.995 -0.165 450.325 0.165 ;
        RECT 448.635 -0.165 448.965 0.165 ;
        RECT 447.275 -0.165 447.605 0.165 ;
        RECT 445.915 -0.165 446.245 0.165 ;
        RECT 444.555 -0.165 444.885 0.165 ;
        RECT 443.195 -0.165 443.525 0.165 ;
        RECT 441.835 -0.165 442.165 0.165 ;
        RECT 440.475 -0.165 440.805 0.165 ;
        RECT 439.115 -0.165 439.445 0.165 ;
        RECT 437.755 -0.165 438.085 0.165 ;
        RECT 436.395 -0.165 436.725 0.165 ;
        RECT 435.035 -0.165 435.365 0.165 ;
        RECT 433.675 -0.165 434.005 0.165 ;
        RECT 432.315 -0.165 432.645 0.165 ;
        RECT 430.955 -0.165 431.285 0.165 ;
        RECT 429.595 -0.165 429.925 0.165 ;
        RECT 428.235 -0.165 428.565 0.165 ;
        RECT 426.875 -0.165 427.205 0.165 ;
        RECT 425.515 -0.165 425.845 0.165 ;
        RECT 424.155 -0.165 424.485 0.165 ;
        RECT 422.795 -0.165 423.125 0.165 ;
        RECT 421.435 -0.165 421.765 0.165 ;
        RECT 420.075 -0.165 420.405 0.165 ;
        RECT 418.715 -0.165 419.045 0.165 ;
        RECT 417.355 -0.165 417.685 0.165 ;
        RECT 415.995 -0.165 416.325 0.165 ;
        RECT 414.635 -0.165 414.965 0.165 ;
        RECT 413.275 -0.165 413.605 0.165 ;
        RECT 411.915 -0.165 412.245 0.165 ;
        RECT 410.555 -0.165 410.885 0.165 ;
        RECT 409.195 -0.165 409.525 0.165 ;
        RECT 407.835 -0.165 408.165 0.165 ;
        RECT 406.475 -0.165 406.805 0.165 ;
        RECT 405.115 -0.165 405.445 0.165 ;
        RECT 403.755 -0.165 404.085 0.165 ;
        RECT 402.395 -0.165 402.725 0.165 ;
        RECT 401.035 -0.165 401.365 0.165 ;
        RECT 399.675 -0.165 400.005 0.165 ;
        RECT 398.315 -0.165 398.645 0.165 ;
        RECT 396.955 -0.165 397.285 0.165 ;
        RECT 395.595 -0.165 395.925 0.165 ;
        RECT 394.235 -0.165 394.565 0.165 ;
        RECT 392.875 -0.165 393.205 0.165 ;
        RECT 391.515 -0.165 391.845 0.165 ;
        RECT 390.155 -0.165 390.485 0.165 ;
        RECT 388.795 -0.165 389.125 0.165 ;
        RECT 387.435 -0.165 387.765 0.165 ;
        RECT 386.075 -0.165 386.405 0.165 ;
        RECT 384.715 -0.165 385.045 0.165 ;
        RECT 383.355 -0.165 383.685 0.165 ;
        RECT 381.995 -0.165 382.325 0.165 ;
        RECT 380.635 -0.165 380.965 0.165 ;
        RECT 379.275 -0.165 379.605 0.165 ;
        RECT 377.915 -0.165 378.245 0.165 ;
        RECT 376.555 -0.165 376.885 0.165 ;
        RECT 375.195 -0.165 375.525 0.165 ;
        RECT 373.835 -0.165 374.165 0.165 ;
        RECT 372.475 -0.165 372.805 0.165 ;
        RECT 371.115 -0.165 371.445 0.165 ;
        RECT 369.755 -0.165 370.085 0.165 ;
        RECT 368.395 -0.165 368.725 0.165 ;
        RECT 367.035 -0.165 367.365 0.165 ;
        RECT 365.675 -0.165 366.005 0.165 ;
        RECT 364.315 -0.165 364.645 0.165 ;
        RECT 362.955 -0.165 363.285 0.165 ;
        RECT 361.595 -0.165 361.925 0.165 ;
        RECT 360.235 -0.165 360.565 0.165 ;
        RECT 358.875 -0.165 359.205 0.165 ;
        RECT 357.515 -0.165 357.845 0.165 ;
        RECT 356.155 -0.165 356.485 0.165 ;
        RECT 354.795 -0.165 355.125 0.165 ;
        RECT 353.435 -0.165 353.765 0.165 ;
        RECT 352.075 -0.165 352.405 0.165 ;
        RECT 350.715 -0.165 351.045 0.165 ;
        RECT 349.355 -0.165 349.685 0.165 ;
        RECT 347.995 -0.165 348.325 0.165 ;
        RECT 346.635 -0.165 346.965 0.165 ;
        RECT 345.275 -0.165 345.605 0.165 ;
        RECT 343.915 -0.165 344.245 0.165 ;
        RECT 342.555 -0.165 342.885 0.165 ;
        RECT 341.195 -0.165 341.525 0.165 ;
        RECT 339.835 -0.165 340.165 0.165 ;
        RECT 338.475 -0.165 338.805 0.165 ;
        RECT 337.115 -0.165 337.445 0.165 ;
        RECT 335.755 -0.165 336.085 0.165 ;
        RECT 334.395 -0.165 334.725 0.165 ;
        RECT 333.035 -0.165 333.365 0.165 ;
        RECT 331.675 -0.165 332.005 0.165 ;
        RECT 330.315 -0.165 330.645 0.165 ;
        RECT 328.955 -0.165 329.285 0.165 ;
        RECT 327.595 -0.165 327.925 0.165 ;
        RECT 326.235 -0.165 326.565 0.165 ;
        RECT 324.875 -0.165 325.205 0.165 ;
        RECT 323.515 -0.165 323.845 0.165 ;
        RECT 322.155 -0.165 322.485 0.165 ;
        RECT 320.795 -0.165 321.125 0.165 ;
        RECT 319.435 -0.165 319.765 0.165 ;
        RECT 318.075 -0.165 318.405 0.165 ;
        RECT 316.715 -0.165 317.045 0.165 ;
        RECT 315.355 -0.165 315.685 0.165 ;
        RECT 313.995 -0.165 314.325 0.165 ;
        RECT 312.635 -0.165 312.965 0.165 ;
        RECT 311.275 -0.165 311.605 0.165 ;
        RECT 309.915 -0.165 310.245 0.165 ;
        RECT 308.555 -0.165 308.885 0.165 ;
        RECT 307.195 -0.165 307.525 0.165 ;
        RECT 305.835 -0.165 306.165 0.165 ;
        RECT 304.475 -0.165 304.805 0.165 ;
        RECT 303.115 -0.165 303.445 0.165 ;
        RECT 301.755 -0.165 302.085 0.165 ;
        RECT 300.395 -0.165 300.725 0.165 ;
        RECT 299.035 -0.165 299.365 0.165 ;
        RECT 297.675 -0.165 298.005 0.165 ;
        RECT 296.315 -0.165 296.645 0.165 ;
        RECT 294.955 -0.165 295.285 0.165 ;
        RECT 293.595 -0.165 293.925 0.165 ;
        RECT 292.235 -0.165 292.565 0.165 ;
        RECT 290.875 -0.165 291.205 0.165 ;
        RECT 289.515 -0.165 289.845 0.165 ;
        RECT 288.155 -0.165 288.485 0.165 ;
        RECT 286.795 -0.165 287.125 0.165 ;
        RECT 285.435 -0.165 285.765 0.165 ;
        RECT 284.075 -0.165 284.405 0.165 ;
        RECT 282.715 -0.165 283.045 0.165 ;
        RECT 281.355 -0.165 281.685 0.165 ;
        RECT 279.995 -0.165 280.325 0.165 ;
        RECT 278.635 -0.165 278.965 0.165 ;
        RECT 277.275 -0.165 277.605 0.165 ;
        RECT 275.915 -0.165 276.245 0.165 ;
        RECT 274.555 -0.165 274.885 0.165 ;
        RECT 273.195 -0.165 273.525 0.165 ;
        RECT 271.835 -0.165 272.165 0.165 ;
        RECT 270.475 -0.165 270.805 0.165 ;
        RECT 269.115 -0.165 269.445 0.165 ;
        RECT 267.755 -0.165 268.085 0.165 ;
        RECT 266.395 -0.165 266.725 0.165 ;
        RECT 265.035 -0.165 265.365 0.165 ;
        RECT 263.675 -0.165 264.005 0.165 ;
        RECT 262.315 -0.165 262.645 0.165 ;
        RECT 260.955 -0.165 261.285 0.165 ;
        RECT 259.595 -0.165 259.925 0.165 ;
        RECT 258.235 -0.165 258.565 0.165 ;
        RECT 256.875 -0.165 257.205 0.165 ;
        RECT 255.515 -0.165 255.845 0.165 ;
        RECT 254.155 -0.165 254.485 0.165 ;
        RECT 252.795 -0.165 253.125 0.165 ;
        RECT 251.435 -0.165 251.765 0.165 ;
        RECT 250.075 -0.165 250.405 0.165 ;
        RECT 248.715 -0.165 249.045 0.165 ;
        RECT 247.355 -0.165 247.685 0.165 ;
        RECT 245.995 -0.165 246.325 0.165 ;
        RECT 244.635 -0.165 244.965 0.165 ;
        RECT 243.275 -0.165 243.605 0.165 ;
        RECT 241.915 -0.165 242.245 0.165 ;
        RECT 240.555 -0.165 240.885 0.165 ;
        RECT 239.195 -0.165 239.525 0.165 ;
        RECT 237.835 -0.165 238.165 0.165 ;
        RECT 236.475 -0.165 236.805 0.165 ;
        RECT 235.115 -0.165 235.445 0.165 ;
        RECT 233.755 -0.165 234.085 0.165 ;
        RECT 232.395 -0.165 232.725 0.165 ;
        RECT 231.035 -0.165 231.365 0.165 ;
        RECT 229.675 -0.165 230.005 0.165 ;
        RECT 228.315 -0.165 228.645 0.165 ;
        RECT 226.955 -0.165 227.285 0.165 ;
        RECT 225.595 -0.165 225.925 0.165 ;
        RECT 224.235 -0.165 224.565 0.165 ;
        RECT 222.875 -0.165 223.205 0.165 ;
        RECT 221.515 -0.165 221.845 0.165 ;
        RECT 220.155 -0.165 220.485 0.165 ;
        RECT 218.795 -0.165 219.125 0.165 ;
        RECT 217.435 -0.165 217.765 0.165 ;
        RECT 216.075 -0.165 216.405 0.165 ;
        RECT 214.715 -0.165 215.045 0.165 ;
        RECT 213.355 -0.165 213.685 0.165 ;
        RECT 211.995 -0.165 212.325 0.165 ;
        RECT 210.635 -0.165 210.965 0.165 ;
        RECT 209.275 -0.165 209.605 0.165 ;
        RECT 207.915 -0.165 208.245 0.165 ;
        RECT 206.555 -0.165 206.885 0.165 ;
        RECT 205.195 -0.165 205.525 0.165 ;
        RECT 203.835 -0.165 204.165 0.165 ;
        RECT 202.475 -0.165 202.805 0.165 ;
        RECT 201.115 -0.165 201.445 0.165 ;
        RECT 199.755 -0.165 200.085 0.165 ;
        RECT 198.395 -0.165 198.725 0.165 ;
        RECT 197.035 -0.165 197.365 0.165 ;
        RECT 195.675 -0.165 196.005 0.165 ;
        RECT 194.315 -0.165 194.645 0.165 ;
        RECT 192.955 -0.165 193.285 0.165 ;
        RECT 191.595 -0.165 191.925 0.165 ;
        RECT 190.235 -0.165 190.565 0.165 ;
        RECT 188.875 -0.165 189.205 0.165 ;
        RECT 187.515 -0.165 187.845 0.165 ;
        RECT 186.155 -0.165 186.485 0.165 ;
        RECT 184.795 -0.165 185.125 0.165 ;
        RECT 183.435 -0.165 183.765 0.165 ;
        RECT 182.075 -0.165 182.405 0.165 ;
        RECT 180.715 -0.165 181.045 0.165 ;
        RECT 179.355 -0.165 179.685 0.165 ;
        RECT 177.995 -0.165 178.325 0.165 ;
        RECT 176.635 -0.165 176.965 0.165 ;
        RECT 175.275 -0.165 175.605 0.165 ;
        RECT 173.915 -0.165 174.245 0.165 ;
        RECT 172.555 -0.165 172.885 0.165 ;
        RECT 171.195 -0.165 171.525 0.165 ;
        RECT 169.835 -0.165 170.165 0.165 ;
        RECT 168.475 -0.165 168.805 0.165 ;
        RECT 167.115 -0.165 167.445 0.165 ;
        RECT 165.755 -0.165 166.085 0.165 ;
        RECT 164.395 -0.165 164.725 0.165 ;
        RECT 163.035 -0.165 163.365 0.165 ;
        RECT 161.675 -0.165 162.005 0.165 ;
        RECT 160.315 -0.165 160.645 0.165 ;
        RECT 158.955 -0.165 159.285 0.165 ;
        RECT 157.595 -0.165 157.925 0.165 ;
        RECT 156.235 -0.165 156.565 0.165 ;
        RECT 154.875 -0.165 155.205 0.165 ;
        RECT 153.515 -0.165 153.845 0.165 ;
        RECT 152.155 -0.165 152.485 0.165 ;
        RECT 150.795 -0.165 151.125 0.165 ;
        RECT 149.435 -0.165 149.765 0.165 ;
        RECT 148.075 -0.165 148.405 0.165 ;
        RECT 146.715 -0.165 147.045 0.165 ;
        RECT 145.355 -0.165 145.685 0.165 ;
        RECT 143.995 -0.165 144.325 0.165 ;
        RECT 142.635 -0.165 142.965 0.165 ;
        RECT 141.275 -0.165 141.605 0.165 ;
        RECT 139.915 -0.165 140.245 0.165 ;
        RECT 138.555 -0.165 138.885 0.165 ;
        RECT 137.195 -0.165 137.525 0.165 ;
        RECT 135.835 -0.165 136.165 0.165 ;
        RECT 134.475 -0.165 134.805 0.165 ;
        RECT 133.115 -0.165 133.445 0.165 ;
        RECT 131.755 -0.165 132.085 0.165 ;
        RECT 130.395 -0.165 130.725 0.165 ;
        RECT 129.035 -0.165 129.365 0.165 ;
        RECT 127.675 -0.165 128.005 0.165 ;
        RECT 126.315 -0.165 126.645 0.165 ;
        RECT 124.955 -0.165 125.285 0.165 ;
        RECT 123.595 -0.165 123.925 0.165 ;
        RECT 122.235 -0.165 122.565 0.165 ;
        RECT 120.875 -0.165 121.205 0.165 ;
        RECT 119.515 -0.165 119.845 0.165 ;
        RECT 118.155 -0.165 118.485 0.165 ;
        RECT 116.795 -0.165 117.125 0.165 ;
        RECT 115.435 -0.165 115.765 0.165 ;
        RECT 114.075 -0.165 114.405 0.165 ;
        RECT 112.715 -0.165 113.045 0.165 ;
        RECT 111.355 -0.165 111.685 0.165 ;
        RECT 109.995 -0.165 110.325 0.165 ;
        RECT 108.635 -0.165 108.965 0.165 ;
        RECT 107.275 -0.165 107.605 0.165 ;
        RECT 105.915 -0.165 106.245 0.165 ;
        RECT 104.555 -0.165 104.885 0.165 ;
        RECT 103.195 -0.165 103.525 0.165 ;
        RECT 101.835 -0.165 102.165 0.165 ;
        RECT 100.475 -0.165 100.805 0.165 ;
        RECT 99.115 -0.165 99.445 0.165 ;
        RECT 97.755 -0.165 98.085 0.165 ;
        RECT 96.395 -0.165 96.725 0.165 ;
        RECT 95.035 -0.165 95.365 0.165 ;
        RECT 93.675 -0.165 94.005 0.165 ;
        RECT 92.315 -0.165 92.645 0.165 ;
        RECT 90.955 -0.165 91.285 0.165 ;
        RECT 89.595 -0.165 89.925 0.165 ;
        RECT 88.235 -0.165 88.565 0.165 ;
        RECT 86.875 -0.165 87.205 0.165 ;
        RECT 85.515 -0.165 85.845 0.165 ;
        RECT 84.155 -0.165 84.485 0.165 ;
        RECT 82.795 -0.165 83.125 0.165 ;
        RECT 81.435 -0.165 81.765 0.165 ;
        RECT 80.075 -0.165 80.405 0.165 ;
        RECT 78.715 -0.165 79.045 0.165 ;
        RECT 77.355 -0.165 77.685 0.165 ;
        RECT 75.995 -0.165 76.325 0.165 ;
        RECT 74.635 -0.165 74.965 0.165 ;
        RECT 73.275 -0.165 73.605 0.165 ;
        RECT 71.915 -0.165 72.245 0.165 ;
        RECT 70.555 -0.165 70.885 0.165 ;
        RECT 69.195 -0.165 69.525 0.165 ;
        RECT 67.835 -0.165 68.165 0.165 ;
        RECT 66.475 -0.165 66.805 0.165 ;
        RECT 65.115 -0.165 65.445 0.165 ;
        RECT 63.755 -0.165 64.085 0.165 ;
        RECT 62.395 -0.165 62.725 0.165 ;
        RECT 61.035 -0.165 61.365 0.165 ;
        RECT 59.675 -0.165 60.005 0.165 ;
        RECT 58.315 -0.165 58.645 0.165 ;
        RECT 56.955 -0.165 57.285 0.165 ;
        RECT 55.595 -0.165 55.925 0.165 ;
        RECT 54.235 -0.165 54.565 0.165 ;
        RECT 52.875 -0.165 53.205 0.165 ;
        RECT 51.515 -0.165 51.845 0.165 ;
        RECT 50.155 -0.165 50.485 0.165 ;
        RECT 48.795 -0.165 49.125 0.165 ;
        RECT 47.435 -0.165 47.765 0.165 ;
        RECT 46.075 -0.165 46.405 0.165 ;
        RECT 44.715 -0.165 45.045 0.165 ;
        RECT 43.355 -0.165 43.685 0.165 ;
        RECT 41.995 -0.165 42.325 0.165 ;
        RECT 40.635 -0.165 40.965 0.165 ;
        RECT 39.275 -0.165 39.605 0.165 ;
        RECT 37.915 -0.165 38.245 0.165 ;
        RECT 36.555 -0.165 36.885 0.165 ;
        RECT 35.195 -0.165 35.525 0.165 ;
        RECT 33.835 -0.165 34.165 0.165 ;
        RECT 32.475 -0.165 32.805 0.165 ;
        RECT 31.115 -0.165 31.445 0.165 ;
        RECT 29.755 -0.165 30.085 0.165 ;
        RECT 28.395 -0.165 28.725 0.165 ;
        RECT 27.035 -0.165 27.365 0.165 ;
        RECT 25.675 -0.165 26.005 0.165 ;
        RECT 24.315 -0.165 24.645 0.165 ;
        RECT 22.955 -0.165 23.285 0.165 ;
        RECT 21.595 -0.165 21.925 0.165 ;
        RECT 20.235 -0.165 20.565 0.165 ;
        RECT 18.875 -0.165 19.205 0.165 ;
        RECT 17.515 -0.165 17.845 0.165 ;
        RECT 16.155 -0.165 16.485 0.165 ;
        RECT 14.795 -0.165 15.125 0.165 ;
        RECT 13.435 -0.165 13.765 0.165 ;
        RECT 12.075 -0.165 12.405 0.165 ;
        RECT 10.715 -0.165 11.045 0.165 ;
        RECT 9.355 -0.165 9.685 0.165 ;
        RECT 7.995 -0.165 8.325 0.165 ;
        RECT 6.635 -0.165 6.965 0.165 ;
        RECT 5.275 -0.165 5.605 0.165 ;
        RECT 3.915 -0.165 4.245 0.165 ;
        RECT 2.555 -0.165 2.885 0.165 ;
        RECT 1.195 -0.165 1.525 0.165 ;
        RECT -0.165 -0.165 0.165 0.165 ;
        RECT -1.525 -0.165 -1.195 0.165 ;
        RECT -1.525 -0.16 678.475 0.16 ;
        RECT 677.115 -0.165 677.445 0.165 ;
        RECT 675.755 -0.165 676.085 0.165 ;
        RECT 674.395 -0.165 674.725 0.165 ;
        RECT 673.035 -0.165 673.365 0.165 ;
        RECT 671.675 -0.165 672.005 0.165 ;
        RECT 670.315 -0.165 670.645 0.165 ;
        RECT 668.955 -0.165 669.285 0.165 ;
        RECT 667.595 -0.165 667.925 0.165 ;
        RECT 666.235 -0.165 666.565 0.165 ;
        RECT 664.875 -0.165 665.205 0.165 ;
        RECT 663.515 -0.165 663.845 0.165 ;
        RECT 662.155 -0.165 662.485 0.165 ;
        RECT 660.795 -0.165 661.125 0.165 ;
        RECT 954.555 -0.165 954.885 0.165 ;
        RECT 678.475 -0.16 954.885 0.16 ;
        RECT 953.195 -0.165 953.525 0.165 ;
        RECT 951.835 -0.165 952.165 0.165 ;
        RECT 950.475 -0.165 950.805 0.165 ;
        RECT 949.115 -0.165 949.445 0.165 ;
        RECT 947.755 -0.165 948.085 0.165 ;
        RECT 946.395 -0.165 946.725 0.165 ;
        RECT 945.035 -0.165 945.365 0.165 ;
        RECT 943.675 -0.165 944.005 0.165 ;
        RECT 942.315 -0.165 942.645 0.165 ;
        RECT 940.955 -0.165 941.285 0.165 ;
        RECT 939.595 -0.165 939.925 0.165 ;
        RECT 938.235 -0.165 938.565 0.165 ;
        RECT 936.875 -0.165 937.205 0.165 ;
        RECT 935.515 -0.165 935.845 0.165 ;
        RECT 934.155 -0.165 934.485 0.165 ;
        RECT 932.795 -0.165 933.125 0.165 ;
        RECT 931.435 -0.165 931.765 0.165 ;
        RECT 930.075 -0.165 930.405 0.165 ;
        RECT 928.715 -0.165 929.045 0.165 ;
        RECT 927.355 -0.165 927.685 0.165 ;
        RECT 925.995 -0.165 926.325 0.165 ;
        RECT 924.635 -0.165 924.965 0.165 ;
        RECT 923.275 -0.165 923.605 0.165 ;
        RECT 921.915 -0.165 922.245 0.165 ;
        RECT 920.555 -0.165 920.885 0.165 ;
        RECT 919.195 -0.165 919.525 0.165 ;
        RECT 917.835 -0.165 918.165 0.165 ;
        RECT 916.475 -0.165 916.805 0.165 ;
        RECT 915.115 -0.165 915.445 0.165 ;
        RECT 913.755 -0.165 914.085 0.165 ;
        RECT 912.395 -0.165 912.725 0.165 ;
        RECT 911.035 -0.165 911.365 0.165 ;
        RECT 909.675 -0.165 910.005 0.165 ;
        RECT 908.315 -0.165 908.645 0.165 ;
        RECT 906.955 -0.165 907.285 0.165 ;
        RECT 905.595 -0.165 905.925 0.165 ;
        RECT 904.235 -0.165 904.565 0.165 ;
        RECT 902.875 -0.165 903.205 0.165 ;
        RECT 901.515 -0.165 901.845 0.165 ;
        RECT 900.155 -0.165 900.485 0.165 ;
        RECT 898.795 -0.165 899.125 0.165 ;
        RECT 897.435 -0.165 897.765 0.165 ;
        RECT 896.075 -0.165 896.405 0.165 ;
        RECT 894.715 -0.165 895.045 0.165 ;
        RECT 893.355 -0.165 893.685 0.165 ;
        RECT 891.995 -0.165 892.325 0.165 ;
        RECT 890.635 -0.165 890.965 0.165 ;
        RECT 889.275 -0.165 889.605 0.165 ;
        RECT 887.915 -0.165 888.245 0.165 ;
        RECT 886.555 -0.165 886.885 0.165 ;
        RECT 885.195 -0.165 885.525 0.165 ;
        RECT 883.835 -0.165 884.165 0.165 ;
        RECT 882.475 -0.165 882.805 0.165 ;
        RECT 881.115 -0.165 881.445 0.165 ;
        RECT 879.755 -0.165 880.085 0.165 ;
        RECT 878.395 -0.165 878.725 0.165 ;
        RECT 877.035 -0.165 877.365 0.165 ;
        RECT 875.675 -0.165 876.005 0.165 ;
        RECT 874.315 -0.165 874.645 0.165 ;
        RECT 872.955 -0.165 873.285 0.165 ;
        RECT 871.595 -0.165 871.925 0.165 ;
        RECT 870.235 -0.165 870.565 0.165 ;
        RECT 868.875 -0.165 869.205 0.165 ;
        RECT 867.515 -0.165 867.845 0.165 ;
        RECT 866.155 -0.165 866.485 0.165 ;
        RECT 864.795 -0.165 865.125 0.165 ;
        RECT 863.435 -0.165 863.765 0.165 ;
        RECT 862.075 -0.165 862.405 0.165 ;
        RECT 860.715 -0.165 861.045 0.165 ;
        RECT 859.355 -0.165 859.685 0.165 ;
        RECT 857.995 -0.165 858.325 0.165 ;
        RECT 856.635 -0.165 856.965 0.165 ;
        RECT 855.275 -0.165 855.605 0.165 ;
        RECT 853.915 -0.165 854.245 0.165 ;
        RECT 852.555 -0.165 852.885 0.165 ;
        RECT 851.195 -0.165 851.525 0.165 ;
        RECT 849.835 -0.165 850.165 0.165 ;
        RECT 848.475 -0.165 848.805 0.165 ;
        RECT 847.115 -0.165 847.445 0.165 ;
        RECT 845.755 -0.165 846.085 0.165 ;
        RECT 844.395 -0.165 844.725 0.165 ;
        RECT 843.035 -0.165 843.365 0.165 ;
        RECT 841.675 -0.165 842.005 0.165 ;
        RECT 840.315 -0.165 840.645 0.165 ;
        RECT 838.955 -0.165 839.285 0.165 ;
        RECT 837.595 -0.165 837.925 0.165 ;
        RECT 836.235 -0.165 836.565 0.165 ;
        RECT 834.875 -0.165 835.205 0.165 ;
        RECT 833.515 -0.165 833.845 0.165 ;
        RECT 832.155 -0.165 832.485 0.165 ;
        RECT 830.795 -0.165 831.125 0.165 ;
        RECT 829.435 -0.165 829.765 0.165 ;
        RECT 828.075 -0.165 828.405 0.165 ;
        RECT 826.715 -0.165 827.045 0.165 ;
        RECT 825.355 -0.165 825.685 0.165 ;
        RECT 823.995 -0.165 824.325 0.165 ;
        RECT 822.635 -0.165 822.965 0.165 ;
        RECT 821.275 -0.165 821.605 0.165 ;
        RECT 819.915 -0.165 820.245 0.165 ;
        RECT 818.555 -0.165 818.885 0.165 ;
        RECT 817.195 -0.165 817.525 0.165 ;
        RECT 815.835 -0.165 816.165 0.165 ;
        RECT 814.475 -0.165 814.805 0.165 ;
        RECT 813.115 -0.165 813.445 0.165 ;
        RECT 811.755 -0.165 812.085 0.165 ;
        RECT 810.395 -0.165 810.725 0.165 ;
        RECT 809.035 -0.165 809.365 0.165 ;
        RECT 807.675 -0.165 808.005 0.165 ;
        RECT 806.315 -0.165 806.645 0.165 ;
        RECT 804.955 -0.165 805.285 0.165 ;
        RECT 803.595 -0.165 803.925 0.165 ;
        RECT 802.235 -0.165 802.565 0.165 ;
        RECT 800.875 -0.165 801.205 0.165 ;
        RECT 799.515 -0.165 799.845 0.165 ;
        RECT 798.155 -0.165 798.485 0.165 ;
        RECT 796.795 -0.165 797.125 0.165 ;
        RECT 795.435 -0.165 795.765 0.165 ;
        RECT 794.075 -0.165 794.405 0.165 ;
        RECT 792.715 -0.165 793.045 0.165 ;
        RECT 791.355 -0.165 791.685 0.165 ;
        RECT 789.995 -0.165 790.325 0.165 ;
        RECT 788.635 -0.165 788.965 0.165 ;
        RECT 787.275 -0.165 787.605 0.165 ;
        RECT 785.915 -0.165 786.245 0.165 ;
        RECT 784.555 -0.165 784.885 0.165 ;
        RECT 783.195 -0.165 783.525 0.165 ;
        RECT 781.835 -0.165 782.165 0.165 ;
        RECT 780.475 -0.165 780.805 0.165 ;
        RECT 779.115 -0.165 779.445 0.165 ;
        RECT 777.755 -0.165 778.085 0.165 ;
        RECT 776.395 -0.165 776.725 0.165 ;
        RECT 775.035 -0.165 775.365 0.165 ;
        RECT 773.675 -0.165 774.005 0.165 ;
        RECT 772.315 -0.165 772.645 0.165 ;
        RECT 770.955 -0.165 771.285 0.165 ;
        RECT 769.595 -0.165 769.925 0.165 ;
        RECT 768.235 -0.165 768.565 0.165 ;
        RECT 766.875 -0.165 767.205 0.165 ;
        RECT 765.515 -0.165 765.845 0.165 ;
        RECT 764.155 -0.165 764.485 0.165 ;
        RECT 762.795 -0.165 763.125 0.165 ;
        RECT 761.435 -0.165 761.765 0.165 ;
        RECT 760.075 -0.165 760.405 0.165 ;
        RECT 758.715 -0.165 759.045 0.165 ;
        RECT 757.355 -0.165 757.685 0.165 ;
        RECT 755.995 -0.165 756.325 0.165 ;
        RECT 754.635 -0.165 754.965 0.165 ;
        RECT 753.275 -0.165 753.605 0.165 ;
        RECT 751.915 -0.165 752.245 0.165 ;
        RECT 750.555 -0.165 750.885 0.165 ;
        RECT 749.195 -0.165 749.525 0.165 ;
        RECT 747.835 -0.165 748.165 0.165 ;
        RECT 746.475 -0.165 746.805 0.165 ;
        RECT 745.115 -0.165 745.445 0.165 ;
        RECT 743.755 -0.165 744.085 0.165 ;
        RECT 742.395 -0.165 742.725 0.165 ;
        RECT 741.035 -0.165 741.365 0.165 ;
        RECT 739.675 -0.165 740.005 0.165 ;
        RECT 738.315 -0.165 738.645 0.165 ;
        RECT 736.955 -0.165 737.285 0.165 ;
        RECT 735.595 -0.165 735.925 0.165 ;
        RECT 734.235 -0.165 734.565 0.165 ;
        RECT 732.875 -0.165 733.205 0.165 ;
        RECT 731.515 -0.165 731.845 0.165 ;
        RECT 730.155 -0.165 730.485 0.165 ;
        RECT 728.795 -0.165 729.125 0.165 ;
        RECT 727.435 -0.165 727.765 0.165 ;
        RECT 726.075 -0.165 726.405 0.165 ;
        RECT 724.715 -0.165 725.045 0.165 ;
        RECT 723.355 -0.165 723.685 0.165 ;
        RECT 721.995 -0.165 722.325 0.165 ;
        RECT 720.635 -0.165 720.965 0.165 ;
        RECT 719.275 -0.165 719.605 0.165 ;
        RECT 717.915 -0.165 718.245 0.165 ;
        RECT 716.555 -0.165 716.885 0.165 ;
        RECT 715.195 -0.165 715.525 0.165 ;
        RECT 713.835 -0.165 714.165 0.165 ;
        RECT 712.475 -0.165 712.805 0.165 ;
        RECT 711.115 -0.165 711.445 0.165 ;
        RECT 709.755 -0.165 710.085 0.165 ;
        RECT 708.395 -0.165 708.725 0.165 ;
        RECT 707.035 -0.165 707.365 0.165 ;
        RECT 705.675 -0.165 706.005 0.165 ;
        RECT 704.315 -0.165 704.645 0.165 ;
        RECT 702.955 -0.165 703.285 0.165 ;
        RECT 701.595 -0.165 701.925 0.165 ;
        RECT 700.235 -0.165 700.565 0.165 ;
        RECT 698.875 -0.165 699.205 0.165 ;
        RECT 697.515 -0.165 697.845 0.165 ;
        RECT 696.155 -0.165 696.485 0.165 ;
        RECT 694.795 -0.165 695.125 0.165 ;
        RECT 693.435 -0.165 693.765 0.165 ;
        RECT 692.075 -0.165 692.405 0.165 ;
        RECT 690.715 -0.165 691.045 0.165 ;
        RECT 689.355 -0.165 689.685 0.165 ;
        RECT 687.995 -0.165 688.325 0.165 ;
        RECT 686.635 -0.165 686.965 0.165 ;
        RECT 685.275 -0.165 685.605 0.165 ;
        RECT 683.915 -0.165 684.245 0.165 ;
        RECT 682.555 -0.165 682.885 0.165 ;
        RECT 681.195 -0.165 681.525 0.165 ;
        RECT 679.835 -0.165 680.165 0.165 ;
        RECT 678.475 -0.165 678.805 0.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.36 -35.52 151.8 -35.2 ;
        RECT 150.795 -35.525 151.125 -35.195 ;
        RECT 149.435 -35.525 149.765 -35.195 ;
        RECT 148.075 -35.525 148.405 -35.195 ;
        RECT 146.715 -35.525 147.045 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.36 -26 155.88 -25.68 ;
        RECT 153.515 -26.005 153.845 -25.675 ;
        RECT 149.435 -26.005 149.765 -25.675 ;
        RECT 148.075 -26.005 148.405 -25.675 ;
        RECT 146.715 -26.005 147.045 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.32 -30.08 166.08 -29.76 ;
        RECT 164.395 -30.085 164.725 -29.755 ;
        RECT 163.035 -30.085 163.365 -29.755 ;
        RECT 161.675 -30.085 162.005 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.56 -23.28 166.76 -22.96 ;
        RECT 164.395 -23.285 164.725 -22.955 ;
        RECT 163.035 -23.285 163.365 -22.955 ;
        RECT 161.675 -23.285 162.005 -22.955 ;
        RECT 160.315 -23.285 160.645 -22.955 ;
        RECT 157.595 -23.285 157.925 -22.955 ;
        RECT 156.235 -23.285 156.565 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.24 -27.36 166.76 -27.04 ;
        RECT 164.395 -27.365 164.725 -27.035 ;
        RECT 163.035 -27.365 163.365 -27.035 ;
        RECT 161.675 -27.365 162.005 -27.035 ;
        RECT 157.595 -27.365 157.925 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.32 -35.52 166.76 -35.2 ;
        RECT 165.755 -35.525 166.085 -35.195 ;
        RECT 164.395 -35.525 164.725 -35.195 ;
        RECT 163.035 -35.525 163.365 -35.195 ;
        RECT 161.675 -35.525 162.005 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.32 -26 170.84 -25.68 ;
        RECT 168.475 -26.005 168.805 -25.675 ;
        RECT 164.395 -26.005 164.725 -25.675 ;
        RECT 163.035 -26.005 163.365 -25.675 ;
        RECT 161.675 -26.005 162.005 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -30.08 181.04 -29.76 ;
        RECT 179.355 -30.085 179.685 -29.755 ;
        RECT 177.995 -30.085 178.325 -29.755 ;
        RECT 176.635 -30.085 176.965 -29.755 ;
        RECT 175.275 -30.085 175.605 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.52 -23.28 181.72 -22.96 ;
        RECT 179.355 -23.285 179.685 -22.955 ;
        RECT 177.995 -23.285 178.325 -22.955 ;
        RECT 176.635 -23.285 176.965 -22.955 ;
        RECT 175.275 -23.285 175.605 -22.955 ;
        RECT 172.555 -23.285 172.885 -22.955 ;
        RECT 171.195 -23.285 171.525 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.2 -27.36 181.72 -27.04 ;
        RECT 179.355 -27.365 179.685 -27.035 ;
        RECT 177.995 -27.365 178.325 -27.035 ;
        RECT 176.635 -27.365 176.965 -27.035 ;
        RECT 175.275 -27.365 175.605 -27.035 ;
        RECT 172.555 -27.365 172.885 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -35.52 181.72 -35.2 ;
        RECT 180.715 -35.525 181.045 -35.195 ;
        RECT 179.355 -35.525 179.685 -35.195 ;
        RECT 177.995 -35.525 178.325 -35.195 ;
        RECT 176.635 -35.525 176.965 -35.195 ;
        RECT 175.275 -35.525 175.605 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -26 185.8 -25.68 ;
        RECT 183.435 -26.005 183.765 -25.675 ;
        RECT 179.355 -26.005 179.685 -25.675 ;
        RECT 177.995 -26.005 178.325 -25.675 ;
        RECT 176.635 -26.005 176.965 -25.675 ;
        RECT 175.275 -26.005 175.605 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.56 -30.08 196 -29.76 ;
        RECT 194.315 -30.085 194.645 -29.755 ;
        RECT 192.955 -30.085 193.285 -29.755 ;
        RECT 191.595 -30.085 191.925 -29.755 ;
        RECT 190.235 -30.085 190.565 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.48 -23.28 196.68 -22.96 ;
        RECT 194.315 -23.285 194.645 -22.955 ;
        RECT 192.955 -23.285 193.285 -22.955 ;
        RECT 191.595 -23.285 191.925 -22.955 ;
        RECT 190.235 -23.285 190.565 -22.955 ;
        RECT 186.155 -23.285 186.485 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.16 -27.36 196.68 -27.04 ;
        RECT 194.315 -27.365 194.645 -27.035 ;
        RECT 192.955 -27.365 193.285 -27.035 ;
        RECT 191.595 -27.365 191.925 -27.035 ;
        RECT 190.235 -27.365 190.565 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.56 -35.52 196.68 -35.2 ;
        RECT 195.675 -35.525 196.005 -35.195 ;
        RECT 194.315 -35.525 194.645 -35.195 ;
        RECT 192.955 -35.525 193.285 -35.195 ;
        RECT 191.595 -35.525 191.925 -35.195 ;
        RECT 190.235 -35.525 190.565 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.56 -26 200.76 -25.68 ;
        RECT 198.395 -26.005 198.725 -25.675 ;
        RECT 194.315 -26.005 194.645 -25.675 ;
        RECT 192.955 -26.005 193.285 -25.675 ;
        RECT 191.595 -26.005 191.925 -25.675 ;
        RECT 190.235 -26.005 190.565 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.52 -30.08 210.96 -29.76 ;
        RECT 209.275 -30.085 209.605 -29.755 ;
        RECT 207.915 -30.085 208.245 -29.755 ;
        RECT 206.555 -30.085 206.885 -29.755 ;
        RECT 205.195 -30.085 205.525 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.44 -23.28 211.64 -22.96 ;
        RECT 209.275 -23.285 209.605 -22.955 ;
        RECT 207.915 -23.285 208.245 -22.955 ;
        RECT 206.555 -23.285 206.885 -22.955 ;
        RECT 205.195 -23.285 205.525 -22.955 ;
        RECT 201.115 -23.285 201.445 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.12 -27.36 211.64 -27.04 ;
        RECT 209.275 -27.365 209.605 -27.035 ;
        RECT 207.915 -27.365 208.245 -27.035 ;
        RECT 206.555 -27.365 206.885 -27.035 ;
        RECT 205.195 -27.365 205.525 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.52 -35.52 211.64 -35.2 ;
        RECT 210.635 -35.525 210.965 -35.195 ;
        RECT 209.275 -35.525 209.605 -35.195 ;
        RECT 207.915 -35.525 208.245 -35.195 ;
        RECT 206.555 -35.525 206.885 -35.195 ;
        RECT 205.195 -35.525 205.525 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.52 -26 215.72 -25.68 ;
        RECT 213.355 -26.005 213.685 -25.675 ;
        RECT 209.275 -26.005 209.605 -25.675 ;
        RECT 207.915 -26.005 208.245 -25.675 ;
        RECT 206.555 -26.005 206.885 -25.675 ;
        RECT 205.195 -26.005 205.525 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.48 -30.08 225.92 -29.76 ;
        RECT 224.235 -30.085 224.565 -29.755 ;
        RECT 222.875 -30.085 223.205 -29.755 ;
        RECT 221.515 -30.085 221.845 -29.755 ;
        RECT 220.155 -30.085 220.485 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.4 -23.28 226.6 -22.96 ;
        RECT 224.235 -23.285 224.565 -22.955 ;
        RECT 222.875 -23.285 223.205 -22.955 ;
        RECT 221.515 -23.285 221.845 -22.955 ;
        RECT 220.155 -23.285 220.485 -22.955 ;
        RECT 216.075 -23.285 216.405 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.08 -27.36 226.6 -27.04 ;
        RECT 224.235 -27.365 224.565 -27.035 ;
        RECT 222.875 -27.365 223.205 -27.035 ;
        RECT 221.515 -27.365 221.845 -27.035 ;
        RECT 220.155 -27.365 220.485 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.48 -35.52 226.6 -35.2 ;
        RECT 225.595 -35.525 225.925 -35.195 ;
        RECT 224.235 -35.525 224.565 -35.195 ;
        RECT 222.875 -35.525 223.205 -35.195 ;
        RECT 221.515 -35.525 221.845 -35.195 ;
        RECT 220.155 -35.525 220.485 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.48 -26 230 -25.68 ;
        RECT 228.315 -26.005 228.645 -25.675 ;
        RECT 224.235 -26.005 224.565 -25.675 ;
        RECT 222.875 -26.005 223.205 -25.675 ;
        RECT 221.515 -26.005 221.845 -25.675 ;
        RECT 220.155 -26.005 220.485 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.44 -30.08 240.88 -29.76 ;
        RECT 239.195 -30.085 239.525 -29.755 ;
        RECT 237.835 -30.085 238.165 -29.755 ;
        RECT 236.475 -30.085 236.805 -29.755 ;
        RECT 235.115 -30.085 235.445 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.36 -23.28 241.56 -22.96 ;
        RECT 239.195 -23.285 239.525 -22.955 ;
        RECT 237.835 -23.285 238.165 -22.955 ;
        RECT 236.475 -23.285 236.805 -22.955 ;
        RECT 235.115 -23.285 235.445 -22.955 ;
        RECT 231.035 -23.285 231.365 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.04 -27.36 241.56 -27.04 ;
        RECT 239.195 -27.365 239.525 -27.035 ;
        RECT 237.835 -27.365 238.165 -27.035 ;
        RECT 236.475 -27.365 236.805 -27.035 ;
        RECT 235.115 -27.365 235.445 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.44 -35.52 241.56 -35.2 ;
        RECT 240.555 -35.525 240.885 -35.195 ;
        RECT 239.195 -35.525 239.525 -35.195 ;
        RECT 237.835 -35.525 238.165 -35.195 ;
        RECT 236.475 -35.525 236.805 -35.195 ;
        RECT 235.115 -35.525 235.445 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.44 -26 244.96 -25.68 ;
        RECT 243.275 -26.005 243.605 -25.675 ;
        RECT 239.195 -26.005 239.525 -25.675 ;
        RECT 237.835 -26.005 238.165 -25.675 ;
        RECT 236.475 -26.005 236.805 -25.675 ;
        RECT 235.115 -26.005 235.445 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -30.08 255.84 -29.76 ;
        RECT 254.155 -30.085 254.485 -29.755 ;
        RECT 252.795 -30.085 253.125 -29.755 ;
        RECT 251.435 -30.085 251.765 -29.755 ;
        RECT 250.075 -30.085 250.405 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.32 -23.28 256.52 -22.96 ;
        RECT 254.155 -23.285 254.485 -22.955 ;
        RECT 252.795 -23.285 253.125 -22.955 ;
        RECT 251.435 -23.285 251.765 -22.955 ;
        RECT 250.075 -23.285 250.405 -22.955 ;
        RECT 245.995 -23.285 246.325 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 246 -27.36 256.52 -27.04 ;
        RECT 254.155 -27.365 254.485 -27.035 ;
        RECT 252.795 -27.365 253.125 -27.035 ;
        RECT 251.435 -27.365 251.765 -27.035 ;
        RECT 250.075 -27.365 250.405 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -35.52 256.52 -35.2 ;
        RECT 255.515 -35.525 255.845 -35.195 ;
        RECT 254.155 -35.525 254.485 -35.195 ;
        RECT 252.795 -35.525 253.125 -35.195 ;
        RECT 251.435 -35.525 251.765 -35.195 ;
        RECT 250.075 -35.525 250.405 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -26 259.92 -25.68 ;
        RECT 258.235 -26.005 258.565 -25.675 ;
        RECT 254.155 -26.005 254.485 -25.675 ;
        RECT 252.795 -26.005 253.125 -25.675 ;
        RECT 251.435 -26.005 251.765 -25.675 ;
        RECT 250.075 -26.005 250.405 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.36 -30.08 270.8 -29.76 ;
        RECT 269.115 -30.085 269.445 -29.755 ;
        RECT 267.755 -30.085 268.085 -29.755 ;
        RECT 266.395 -30.085 266.725 -29.755 ;
        RECT 265.035 -30.085 265.365 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.28 -23.28 271.48 -22.96 ;
        RECT 269.115 -23.285 269.445 -22.955 ;
        RECT 267.755 -23.285 268.085 -22.955 ;
        RECT 266.395 -23.285 266.725 -22.955 ;
        RECT 265.035 -23.285 265.365 -22.955 ;
        RECT 260.955 -23.285 261.285 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.28 -27.36 271.48 -27.04 ;
        RECT 269.115 -27.365 269.445 -27.035 ;
        RECT 267.755 -27.365 268.085 -27.035 ;
        RECT 266.395 -27.365 266.725 -27.035 ;
        RECT 265.035 -27.365 265.365 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.36 -35.52 271.48 -35.2 ;
        RECT 270.475 -35.525 270.805 -35.195 ;
        RECT 269.115 -35.525 269.445 -35.195 ;
        RECT 267.755 -35.525 268.085 -35.195 ;
        RECT 266.395 -35.525 266.725 -35.195 ;
        RECT 265.035 -35.525 265.365 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.36 -26 274.88 -25.68 ;
        RECT 273.195 -26.005 273.525 -25.675 ;
        RECT 269.115 -26.005 269.445 -25.675 ;
        RECT 267.755 -26.005 268.085 -25.675 ;
        RECT 266.395 -26.005 266.725 -25.675 ;
        RECT 265.035 -26.005 265.365 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.32 -30.08 285.76 -29.76 ;
        RECT 284.075 -30.085 284.405 -29.755 ;
        RECT 282.715 -30.085 283.045 -29.755 ;
        RECT 281.355 -30.085 281.685 -29.755 ;
        RECT 279.995 -30.085 280.325 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.56 -23.28 286.44 -22.96 ;
        RECT 284.075 -23.285 284.405 -22.955 ;
        RECT 282.715 -23.285 283.045 -22.955 ;
        RECT 281.355 -23.285 281.685 -22.955 ;
        RECT 279.995 -23.285 280.325 -22.955 ;
        RECT 275.915 -23.285 276.245 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.24 -27.36 286.44 -27.04 ;
        RECT 284.075 -27.365 284.405 -27.035 ;
        RECT 282.715 -27.365 283.045 -27.035 ;
        RECT 281.355 -27.365 281.685 -27.035 ;
        RECT 279.995 -27.365 280.325 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.32 -35.52 286.44 -35.2 ;
        RECT 285.435 -35.525 285.765 -35.195 ;
        RECT 284.075 -35.525 284.405 -35.195 ;
        RECT 282.715 -35.525 283.045 -35.195 ;
        RECT 281.355 -35.525 281.685 -35.195 ;
        RECT 279.995 -35.525 280.325 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.32 -26 289.84 -25.68 ;
        RECT 288.155 -26.005 288.485 -25.675 ;
        RECT 284.075 -26.005 284.405 -25.675 ;
        RECT 282.715 -26.005 283.045 -25.675 ;
        RECT 281.355 -26.005 281.685 -25.675 ;
        RECT 279.995 -26.005 280.325 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.52 -23.28 300.72 -22.96 ;
        RECT 299.035 -23.285 299.365 -22.955 ;
        RECT 297.675 -23.285 298.005 -22.955 ;
        RECT 296.315 -23.285 296.645 -22.955 ;
        RECT 294.955 -23.285 295.285 -22.955 ;
        RECT 290.875 -23.285 291.205 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -27.36 300.72 -27.04 ;
        RECT 299.035 -27.365 299.365 -27.035 ;
        RECT 297.675 -27.365 298.005 -27.035 ;
        RECT 296.315 -27.365 296.645 -27.035 ;
        RECT 294.955 -27.365 295.285 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.28 -30.08 300.72 -29.76 ;
        RECT 299.035 -30.085 299.365 -29.755 ;
        RECT 297.675 -30.085 298.005 -29.755 ;
        RECT 296.315 -30.085 296.645 -29.755 ;
        RECT 294.955 -30.085 295.285 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 -35.525 300.725 -35.195 ;
        RECT 294.28 -35.52 300.725 -35.2 ;
        RECT 299.035 -35.525 299.365 -35.195 ;
        RECT 297.675 -35.525 298.005 -35.195 ;
        RECT 296.315 -35.525 296.645 -35.195 ;
        RECT 294.955 -35.525 295.285 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.28 -26 304.8 -25.68 ;
        RECT 303.115 -26.005 303.445 -25.675 ;
        RECT 299.035 -26.005 299.365 -25.675 ;
        RECT 297.675 -26.005 298.005 -25.675 ;
        RECT 296.315 -26.005 296.645 -25.675 ;
        RECT 294.955 -26.005 295.285 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.24 -30.08 315 -29.76 ;
        RECT 313.995 -30.085 314.325 -29.755 ;
        RECT 312.635 -30.085 312.965 -29.755 ;
        RECT 311.275 -30.085 311.605 -29.755 ;
        RECT 309.915 -30.085 310.245 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.48 -23.28 315.68 -22.96 ;
        RECT 313.995 -23.285 314.325 -22.955 ;
        RECT 312.635 -23.285 312.965 -22.955 ;
        RECT 311.275 -23.285 311.605 -22.955 ;
        RECT 309.915 -23.285 310.245 -22.955 ;
        RECT 305.835 -23.285 306.165 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.16 -27.36 315.68 -27.04 ;
        RECT 313.995 -27.365 314.325 -27.035 ;
        RECT 312.635 -27.365 312.965 -27.035 ;
        RECT 311.275 -27.365 311.605 -27.035 ;
        RECT 309.915 -27.365 310.245 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 -35.525 315.685 -35.195 ;
        RECT 309.24 -35.52 315.685 -35.2 ;
        RECT 313.995 -35.525 314.325 -35.195 ;
        RECT 312.635 -35.525 312.965 -35.195 ;
        RECT 311.275 -35.525 311.605 -35.195 ;
        RECT 309.915 -35.525 310.245 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.24 -26 319.76 -25.68 ;
        RECT 318.075 -26.005 318.405 -25.675 ;
        RECT 316.715 -26.005 317.045 -25.675 ;
        RECT 313.995 -26.005 314.325 -25.675 ;
        RECT 312.635 -26.005 312.965 -25.675 ;
        RECT 311.275 -26.005 311.605 -25.675 ;
        RECT 309.915 -26.005 310.245 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.2 -30.08 329.96 -29.76 ;
        RECT 328.955 -30.085 329.285 -29.755 ;
        RECT 327.595 -30.085 327.925 -29.755 ;
        RECT 326.235 -30.085 326.565 -29.755 ;
        RECT 324.875 -30.085 325.205 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.44 -23.28 330.64 -22.96 ;
        RECT 328.955 -23.285 329.285 -22.955 ;
        RECT 327.595 -23.285 327.925 -22.955 ;
        RECT 326.235 -23.285 326.565 -22.955 ;
        RECT 324.875 -23.285 325.205 -22.955 ;
        RECT 320.795 -23.285 321.125 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.12 -27.36 330.64 -27.04 ;
        RECT 328.955 -27.365 329.285 -27.035 ;
        RECT 327.595 -27.365 327.925 -27.035 ;
        RECT 326.235 -27.365 326.565 -27.035 ;
        RECT 324.875 -27.365 325.205 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 -35.525 330.645 -35.195 ;
        RECT 324.2 -35.52 330.645 -35.2 ;
        RECT 328.955 -35.525 329.285 -35.195 ;
        RECT 327.595 -35.525 327.925 -35.195 ;
        RECT 326.235 -35.525 326.565 -35.195 ;
        RECT 324.875 -35.525 325.205 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.2 -26 334.72 -25.68 ;
        RECT 333.035 -26.005 333.365 -25.675 ;
        RECT 331.675 -26.005 332.005 -25.675 ;
        RECT 328.955 -26.005 329.285 -25.675 ;
        RECT 327.595 -26.005 327.925 -25.675 ;
        RECT 326.235 -26.005 326.565 -25.675 ;
        RECT 324.875 -26.005 325.205 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.16 -30.08 344.92 -29.76 ;
        RECT 343.915 -30.085 344.245 -29.755 ;
        RECT 342.555 -30.085 342.885 -29.755 ;
        RECT 341.195 -30.085 341.525 -29.755 ;
        RECT 339.835 -30.085 340.165 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.4 -23.28 345.6 -22.96 ;
        RECT 343.915 -23.285 344.245 -22.955 ;
        RECT 342.555 -23.285 342.885 -22.955 ;
        RECT 341.195 -23.285 341.525 -22.955 ;
        RECT 339.835 -23.285 340.165 -22.955 ;
        RECT 335.755 -23.285 336.085 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.08 -27.36 345.6 -27.04 ;
        RECT 343.915 -27.365 344.245 -27.035 ;
        RECT 342.555 -27.365 342.885 -27.035 ;
        RECT 341.195 -27.365 341.525 -27.035 ;
        RECT 339.835 -27.365 340.165 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 -35.525 345.605 -35.195 ;
        RECT 339.16 -35.52 345.605 -35.2 ;
        RECT 343.915 -35.525 344.245 -35.195 ;
        RECT 342.555 -35.525 342.885 -35.195 ;
        RECT 341.195 -35.525 341.525 -35.195 ;
        RECT 339.835 -35.525 340.165 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.16 -26 349.68 -25.68 ;
        RECT 347.995 -26.005 348.325 -25.675 ;
        RECT 346.635 -26.005 346.965 -25.675 ;
        RECT 343.915 -26.005 344.245 -25.675 ;
        RECT 342.555 -26.005 342.885 -25.675 ;
        RECT 341.195 -26.005 341.525 -25.675 ;
        RECT 339.835 -26.005 340.165 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.44 -30.08 359.88 -29.76 ;
        RECT 358.875 -30.085 359.205 -29.755 ;
        RECT 357.515 -30.085 357.845 -29.755 ;
        RECT 356.155 -30.085 356.485 -29.755 ;
        RECT 354.795 -30.085 355.125 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.36 -23.28 360.56 -22.96 ;
        RECT 358.875 -23.285 359.205 -22.955 ;
        RECT 357.515 -23.285 357.845 -22.955 ;
        RECT 356.155 -23.285 356.485 -22.955 ;
        RECT 354.795 -23.285 355.125 -22.955 ;
        RECT 353.435 -23.285 353.765 -22.955 ;
        RECT 350.715 -23.285 351.045 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.04 -27.36 360.56 -27.04 ;
        RECT 358.875 -27.365 359.205 -27.035 ;
        RECT 357.515 -27.365 357.845 -27.035 ;
        RECT 356.155 -27.365 356.485 -27.035 ;
        RECT 354.795 -27.365 355.125 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 -35.525 360.565 -35.195 ;
        RECT 353.44 -35.52 360.565 -35.2 ;
        RECT 358.875 -35.525 359.205 -35.195 ;
        RECT 357.515 -35.525 357.845 -35.195 ;
        RECT 356.155 -35.525 356.485 -35.195 ;
        RECT 354.795 -35.525 355.125 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.44 -26 364.64 -25.68 ;
        RECT 362.955 -26.005 363.285 -25.675 ;
        RECT 361.595 -26.005 361.925 -25.675 ;
        RECT 358.875 -26.005 359.205 -25.675 ;
        RECT 357.515 -26.005 357.845 -25.675 ;
        RECT 356.155 -26.005 356.485 -25.675 ;
        RECT 354.795 -26.005 355.125 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.4 -30.08 374.84 -29.76 ;
        RECT 373.835 -30.085 374.165 -29.755 ;
        RECT 372.475 -30.085 372.805 -29.755 ;
        RECT 371.115 -30.085 371.445 -29.755 ;
        RECT 369.755 -30.085 370.085 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.32 -23.28 375.52 -22.96 ;
        RECT 373.835 -23.285 374.165 -22.955 ;
        RECT 372.475 -23.285 372.805 -22.955 ;
        RECT 371.115 -23.285 371.445 -22.955 ;
        RECT 369.755 -23.285 370.085 -22.955 ;
        RECT 368.395 -23.285 368.725 -22.955 ;
        RECT 365.675 -23.285 366.005 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 365 -27.36 375.52 -27.04 ;
        RECT 373.835 -27.365 374.165 -27.035 ;
        RECT 372.475 -27.365 372.805 -27.035 ;
        RECT 371.115 -27.365 371.445 -27.035 ;
        RECT 369.755 -27.365 370.085 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.195 -35.525 375.525 -35.195 ;
        RECT 368.4 -35.52 375.525 -35.2 ;
        RECT 373.835 -35.525 374.165 -35.195 ;
        RECT 372.475 -35.525 372.805 -35.195 ;
        RECT 371.115 -35.525 371.445 -35.195 ;
        RECT 369.755 -35.525 370.085 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.4 -26 379.6 -25.68 ;
        RECT 377.915 -26.005 378.245 -25.675 ;
        RECT 376.555 -26.005 376.885 -25.675 ;
        RECT 373.835 -26.005 374.165 -25.675 ;
        RECT 372.475 -26.005 372.805 -25.675 ;
        RECT 371.115 -26.005 371.445 -25.675 ;
        RECT 369.755 -26.005 370.085 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.36 -30.08 389.8 -29.76 ;
        RECT 388.795 -30.085 389.125 -29.755 ;
        RECT 387.435 -30.085 387.765 -29.755 ;
        RECT 386.075 -30.085 386.405 -29.755 ;
        RECT 384.715 -30.085 385.045 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.28 -23.28 390.48 -22.96 ;
        RECT 388.795 -23.285 389.125 -22.955 ;
        RECT 387.435 -23.285 387.765 -22.955 ;
        RECT 386.075 -23.285 386.405 -22.955 ;
        RECT 384.715 -23.285 385.045 -22.955 ;
        RECT 383.355 -23.285 383.685 -22.955 ;
        RECT 380.635 -23.285 380.965 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.96 -27.36 390.48 -27.04 ;
        RECT 388.795 -27.365 389.125 -27.035 ;
        RECT 387.435 -27.365 387.765 -27.035 ;
        RECT 386.075 -27.365 386.405 -27.035 ;
        RECT 384.715 -27.365 385.045 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.155 -35.525 390.485 -35.195 ;
        RECT 383.36 -35.52 390.485 -35.2 ;
        RECT 388.795 -35.525 389.125 -35.195 ;
        RECT 387.435 -35.525 387.765 -35.195 ;
        RECT 386.075 -35.525 386.405 -35.195 ;
        RECT 384.715 -35.525 385.045 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.36 -26 393.88 -25.68 ;
        RECT 392.875 -26.005 393.205 -25.675 ;
        RECT 391.515 -26.005 391.845 -25.675 ;
        RECT 388.795 -26.005 389.125 -25.675 ;
        RECT 387.435 -26.005 387.765 -25.675 ;
        RECT 386.075 -26.005 386.405 -25.675 ;
        RECT 384.715 -26.005 385.045 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.32 -30.08 404.76 -29.76 ;
        RECT 403.755 -30.085 404.085 -29.755 ;
        RECT 402.395 -30.085 402.725 -29.755 ;
        RECT 401.035 -30.085 401.365 -29.755 ;
        RECT 399.675 -30.085 400.005 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.24 -23.28 405.44 -22.96 ;
        RECT 403.755 -23.285 404.085 -22.955 ;
        RECT 402.395 -23.285 402.725 -22.955 ;
        RECT 401.035 -23.285 401.365 -22.955 ;
        RECT 399.675 -23.285 400.005 -22.955 ;
        RECT 398.315 -23.285 398.645 -22.955 ;
        RECT 395.595 -23.285 395.925 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.92 -27.36 405.44 -27.04 ;
        RECT 403.755 -27.365 404.085 -27.035 ;
        RECT 402.395 -27.365 402.725 -27.035 ;
        RECT 401.035 -27.365 401.365 -27.035 ;
        RECT 399.675 -27.365 400.005 -27.035 ;
        RECT 395.595 -27.365 395.925 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 405.115 -35.525 405.445 -35.195 ;
        RECT 398.32 -35.52 405.445 -35.2 ;
        RECT 403.755 -35.525 404.085 -35.195 ;
        RECT 402.395 -35.525 402.725 -35.195 ;
        RECT 401.035 -35.525 401.365 -35.195 ;
        RECT 399.675 -35.525 400.005 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 398.32 -26 408.84 -25.68 ;
        RECT 407.835 -26.005 408.165 -25.675 ;
        RECT 406.475 -26.005 406.805 -25.675 ;
        RECT 403.755 -26.005 404.085 -25.675 ;
        RECT 402.395 -26.005 402.725 -25.675 ;
        RECT 401.035 -26.005 401.365 -25.675 ;
        RECT 399.675 -26.005 400.005 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.28 -30.08 419.72 -29.76 ;
        RECT 418.715 -30.085 419.045 -29.755 ;
        RECT 417.355 -30.085 417.685 -29.755 ;
        RECT 415.995 -30.085 416.325 -29.755 ;
        RECT 414.635 -30.085 414.965 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.2 -23.28 420.4 -22.96 ;
        RECT 418.715 -23.285 419.045 -22.955 ;
        RECT 417.355 -23.285 417.685 -22.955 ;
        RECT 415.995 -23.285 416.325 -22.955 ;
        RECT 414.635 -23.285 414.965 -22.955 ;
        RECT 413.275 -23.285 413.605 -22.955 ;
        RECT 410.555 -23.285 410.885 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 409.88 -27.36 420.4 -27.04 ;
        RECT 418.715 -27.365 419.045 -27.035 ;
        RECT 417.355 -27.365 417.685 -27.035 ;
        RECT 415.995 -27.365 416.325 -27.035 ;
        RECT 414.635 -27.365 414.965 -27.035 ;
        RECT 410.555 -27.365 410.885 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 420.075 -35.525 420.405 -35.195 ;
        RECT 413.28 -35.52 420.405 -35.2 ;
        RECT 418.715 -35.525 419.045 -35.195 ;
        RECT 417.355 -35.525 417.685 -35.195 ;
        RECT 415.995 -35.525 416.325 -35.195 ;
        RECT 414.635 -35.525 414.965 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 413.28 -26 423.8 -25.68 ;
        RECT 421.435 -26.005 421.765 -25.675 ;
        RECT 418.715 -26.005 419.045 -25.675 ;
        RECT 417.355 -26.005 417.685 -25.675 ;
        RECT 415.995 -26.005 416.325 -25.675 ;
        RECT 414.635 -26.005 414.965 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.24 -30.08 434.68 -29.76 ;
        RECT 433.675 -30.085 434.005 -29.755 ;
        RECT 432.315 -30.085 432.645 -29.755 ;
        RECT 430.955 -30.085 431.285 -29.755 ;
        RECT 429.595 -30.085 429.925 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.155 -23.28 435.36 -22.96 ;
        RECT 433.675 -23.285 434.005 -22.955 ;
        RECT 432.315 -23.285 432.645 -22.955 ;
        RECT 430.955 -23.285 431.285 -22.955 ;
        RECT 429.595 -23.285 429.925 -22.955 ;
        RECT 428.235 -23.285 428.565 -22.955 ;
        RECT 425.515 -23.285 425.845 -22.955 ;
        RECT 424.155 -23.285 424.485 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 424.16 -27.36 435.36 -27.04 ;
        RECT 433.675 -27.365 434.005 -27.035 ;
        RECT 432.315 -27.365 432.645 -27.035 ;
        RECT 430.955 -27.365 431.285 -27.035 ;
        RECT 429.595 -27.365 429.925 -27.035 ;
        RECT 425.515 -27.365 425.845 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 435.035 -35.525 435.365 -35.195 ;
        RECT 428.24 -35.52 435.365 -35.2 ;
        RECT 433.675 -35.525 434.005 -35.195 ;
        RECT 432.315 -35.525 432.645 -35.195 ;
        RECT 430.955 -35.525 431.285 -35.195 ;
        RECT 429.595 -35.525 429.925 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 428.24 -26 438.76 -25.68 ;
        RECT 436.395 -26.005 436.725 -25.675 ;
        RECT 433.675 -26.005 434.005 -25.675 ;
        RECT 432.315 -26.005 432.645 -25.675 ;
        RECT 430.955 -26.005 431.285 -25.675 ;
        RECT 429.595 -26.005 429.925 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.2 -30.08 449.64 -29.76 ;
        RECT 448.635 -30.085 448.965 -29.755 ;
        RECT 447.275 -30.085 447.605 -29.755 ;
        RECT 445.915 -30.085 446.245 -29.755 ;
        RECT 444.555 -30.085 444.885 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 438.44 -23.28 450.32 -22.96 ;
        RECT 448.635 -23.285 448.965 -22.955 ;
        RECT 447.275 -23.285 447.605 -22.955 ;
        RECT 445.915 -23.285 446.245 -22.955 ;
        RECT 444.555 -23.285 444.885 -22.955 ;
        RECT 443.195 -23.285 443.525 -22.955 ;
        RECT 440.475 -23.285 440.805 -22.955 ;
        RECT 439.115 -23.285 439.445 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 439.12 -27.36 450.32 -27.04 ;
        RECT 448.635 -27.365 448.965 -27.035 ;
        RECT 447.275 -27.365 447.605 -27.035 ;
        RECT 445.915 -27.365 446.245 -27.035 ;
        RECT 444.555 -27.365 444.885 -27.035 ;
        RECT 440.475 -27.365 440.805 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 449.995 -35.525 450.325 -35.195 ;
        RECT 443.2 -35.52 450.325 -35.2 ;
        RECT 448.635 -35.525 448.965 -35.195 ;
        RECT 447.275 -35.525 447.605 -35.195 ;
        RECT 445.915 -35.525 446.245 -35.195 ;
        RECT 444.555 -35.525 444.885 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 443.2 -26 453.72 -25.68 ;
        RECT 451.355 -26.005 451.685 -25.675 ;
        RECT 448.635 -26.005 448.965 -25.675 ;
        RECT 447.275 -26.005 447.605 -25.675 ;
        RECT 445.915 -26.005 446.245 -25.675 ;
        RECT 444.555 -26.005 444.885 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 453.4 -23.28 464.6 -22.96 ;
        RECT 463.595 -23.285 463.925 -22.955 ;
        RECT 462.235 -23.285 462.565 -22.955 ;
        RECT 460.875 -23.285 461.205 -22.955 ;
        RECT 459.515 -23.285 459.845 -22.955 ;
        RECT 458.155 -23.285 458.485 -22.955 ;
        RECT 455.435 -23.285 455.765 -22.955 ;
        RECT 454.075 -23.285 454.405 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 454.08 -27.36 464.6 -27.04 ;
        RECT 463.595 -27.365 463.925 -27.035 ;
        RECT 462.235 -27.365 462.565 -27.035 ;
        RECT 460.875 -27.365 461.205 -27.035 ;
        RECT 459.515 -27.365 459.845 -27.035 ;
        RECT 455.435 -27.365 455.765 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.16 -30.08 464.6 -29.76 ;
        RECT 463.595 -30.085 463.925 -29.755 ;
        RECT 462.235 -30.085 462.565 -29.755 ;
        RECT 460.875 -30.085 461.205 -29.755 ;
        RECT 459.515 -30.085 459.845 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.16 -35.52 464.6 -35.2 ;
        RECT 463.595 -35.525 463.925 -35.195 ;
        RECT 462.235 -35.525 462.565 -35.195 ;
        RECT 460.875 -35.525 461.205 -35.195 ;
        RECT 459.515 -35.525 459.845 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 458.16 -26 468.68 -25.68 ;
        RECT 466.315 -26.005 466.645 -25.675 ;
        RECT 463.595 -26.005 463.925 -25.675 ;
        RECT 462.235 -26.005 462.565 -25.675 ;
        RECT 460.875 -26.005 461.205 -25.675 ;
        RECT 459.515 -26.005 459.845 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.12 -30.08 478.88 -29.76 ;
        RECT 477.195 -30.085 477.525 -29.755 ;
        RECT 475.835 -30.085 476.165 -29.755 ;
        RECT 474.475 -30.085 474.805 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 468.36 -23.28 479.56 -22.96 ;
        RECT 477.195 -23.285 477.525 -22.955 ;
        RECT 475.835 -23.285 476.165 -22.955 ;
        RECT 474.475 -23.285 474.805 -22.955 ;
        RECT 473.115 -23.285 473.445 -22.955 ;
        RECT 470.395 -23.285 470.725 -22.955 ;
        RECT 469.035 -23.285 469.365 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 469.04 -27.36 479.56 -27.04 ;
        RECT 477.195 -27.365 477.525 -27.035 ;
        RECT 475.835 -27.365 476.165 -27.035 ;
        RECT 474.475 -27.365 474.805 -27.035 ;
        RECT 470.395 -27.365 470.725 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.12 -35.52 479.56 -35.2 ;
        RECT 478.555 -35.525 478.885 -35.195 ;
        RECT 477.195 -35.525 477.525 -35.195 ;
        RECT 475.835 -35.525 476.165 -35.195 ;
        RECT 474.475 -35.525 474.805 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 473.12 -26 483.64 -25.68 ;
        RECT 481.275 -26.005 481.605 -25.675 ;
        RECT 477.195 -26.005 477.525 -25.675 ;
        RECT 475.835 -26.005 476.165 -25.675 ;
        RECT 474.475 -26.005 474.805 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.08 -30.08 493.84 -29.76 ;
        RECT 492.155 -30.085 492.485 -29.755 ;
        RECT 490.795 -30.085 491.125 -29.755 ;
        RECT 489.435 -30.085 489.765 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 483.32 -23.28 494.52 -22.96 ;
        RECT 492.155 -23.285 492.485 -22.955 ;
        RECT 490.795 -23.285 491.125 -22.955 ;
        RECT 489.435 -23.285 489.765 -22.955 ;
        RECT 488.075 -23.285 488.405 -22.955 ;
        RECT 485.355 -23.285 485.685 -22.955 ;
        RECT 483.995 -23.285 484.325 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 484 -27.36 494.52 -27.04 ;
        RECT 492.155 -27.365 492.485 -27.035 ;
        RECT 490.795 -27.365 491.125 -27.035 ;
        RECT 489.435 -27.365 489.765 -27.035 ;
        RECT 485.355 -27.365 485.685 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.08 -35.52 494.52 -35.2 ;
        RECT 493.515 -35.525 493.845 -35.195 ;
        RECT 492.155 -35.525 492.485 -35.195 ;
        RECT 490.795 -35.525 491.125 -35.195 ;
        RECT 489.435 -35.525 489.765 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 488.08 -26 498.6 -25.68 ;
        RECT 496.235 -26.005 496.565 -25.675 ;
        RECT 492.155 -26.005 492.485 -25.675 ;
        RECT 490.795 -26.005 491.125 -25.675 ;
        RECT 489.435 -26.005 489.765 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.04 -30.08 508.8 -29.76 ;
        RECT 507.115 -30.085 507.445 -29.755 ;
        RECT 505.755 -30.085 506.085 -29.755 ;
        RECT 504.395 -30.085 504.725 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.28 -23.28 509.48 -22.96 ;
        RECT 507.115 -23.285 507.445 -22.955 ;
        RECT 505.755 -23.285 506.085 -22.955 ;
        RECT 504.395 -23.285 504.725 -22.955 ;
        RECT 503.035 -23.285 503.365 -22.955 ;
        RECT 500.315 -23.285 500.645 -22.955 ;
        RECT 498.955 -23.285 499.285 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 498.96 -27.36 509.48 -27.04 ;
        RECT 507.115 -27.365 507.445 -27.035 ;
        RECT 505.755 -27.365 506.085 -27.035 ;
        RECT 504.395 -27.365 504.725 -27.035 ;
        RECT 500.315 -27.365 500.645 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.04 -35.52 509.48 -35.2 ;
        RECT 508.475 -35.525 508.805 -35.195 ;
        RECT 507.115 -35.525 507.445 -35.195 ;
        RECT 505.755 -35.525 506.085 -35.195 ;
        RECT 504.395 -35.525 504.725 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 503.04 -26 513.56 -25.68 ;
        RECT 511.195 -26.005 511.525 -25.675 ;
        RECT 507.115 -26.005 507.445 -25.675 ;
        RECT 505.755 -26.005 506.085 -25.675 ;
        RECT 504.395 -26.005 504.725 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.995 -30.08 523.76 -29.76 ;
        RECT 522.075 -30.085 522.405 -29.755 ;
        RECT 520.715 -30.085 521.045 -29.755 ;
        RECT 519.355 -30.085 519.685 -29.755 ;
        RECT 517.995 -30.085 518.325 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.24 -23.28 524.44 -22.96 ;
        RECT 522.075 -23.285 522.405 -22.955 ;
        RECT 520.715 -23.285 521.045 -22.955 ;
        RECT 519.355 -23.285 519.685 -22.955 ;
        RECT 517.995 -23.285 518.325 -22.955 ;
        RECT 515.275 -23.285 515.605 -22.955 ;
        RECT 513.915 -23.285 514.245 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 513.92 -27.36 524.44 -27.04 ;
        RECT 522.075 -27.365 522.405 -27.035 ;
        RECT 520.715 -27.365 521.045 -27.035 ;
        RECT 519.355 -27.365 519.685 -27.035 ;
        RECT 517.995 -27.365 518.325 -27.035 ;
        RECT 515.275 -27.365 515.605 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.995 -35.52 524.44 -35.2 ;
        RECT 523.435 -35.525 523.765 -35.195 ;
        RECT 522.075 -35.525 522.405 -35.195 ;
        RECT 520.715 -35.525 521.045 -35.195 ;
        RECT 519.355 -35.525 519.685 -35.195 ;
        RECT 517.995 -35.525 518.325 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 517.995 -26 528.52 -25.68 ;
        RECT 526.155 -26.005 526.485 -25.675 ;
        RECT 522.075 -26.005 522.405 -25.675 ;
        RECT 520.715 -26.005 521.045 -25.675 ;
        RECT 519.355 -26.005 519.685 -25.675 ;
        RECT 517.995 -26.005 518.325 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.28 -30.08 538.72 -29.76 ;
        RECT 537.035 -30.085 537.365 -29.755 ;
        RECT 535.675 -30.085 536.005 -29.755 ;
        RECT 534.315 -30.085 534.645 -29.755 ;
        RECT 532.955 -30.085 533.285 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.2 -23.28 539.4 -22.96 ;
        RECT 537.035 -23.285 537.365 -22.955 ;
        RECT 535.675 -23.285 536.005 -22.955 ;
        RECT 534.315 -23.285 534.645 -22.955 ;
        RECT 532.955 -23.285 533.285 -22.955 ;
        RECT 528.875 -23.285 529.205 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 528.88 -27.36 539.4 -27.04 ;
        RECT 537.035 -27.365 537.365 -27.035 ;
        RECT 535.675 -27.365 536.005 -27.035 ;
        RECT 534.315 -27.365 534.645 -27.035 ;
        RECT 532.955 -27.365 533.285 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.28 -35.52 539.4 -35.2 ;
        RECT 538.395 -35.525 538.725 -35.195 ;
        RECT 537.035 -35.525 537.365 -35.195 ;
        RECT 535.675 -35.525 536.005 -35.195 ;
        RECT 534.315 -35.525 534.645 -35.195 ;
        RECT 532.955 -35.525 533.285 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 532.28 -26 543.48 -25.68 ;
        RECT 541.115 -26.005 541.445 -25.675 ;
        RECT 537.035 -26.005 537.365 -25.675 ;
        RECT 535.675 -26.005 536.005 -25.675 ;
        RECT 534.315 -26.005 534.645 -25.675 ;
        RECT 532.955 -26.005 533.285 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.24 -30.08 553.68 -29.76 ;
        RECT 551.995 -30.085 552.325 -29.755 ;
        RECT 550.635 -30.085 550.965 -29.755 ;
        RECT 549.275 -30.085 549.605 -29.755 ;
        RECT 547.915 -30.085 548.245 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.16 -23.28 554.36 -22.96 ;
        RECT 551.995 -23.285 552.325 -22.955 ;
        RECT 550.635 -23.285 550.965 -22.955 ;
        RECT 549.275 -23.285 549.605 -22.955 ;
        RECT 547.915 -23.285 548.245 -22.955 ;
        RECT 543.835 -23.285 544.165 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 543.84 -27.36 554.36 -27.04 ;
        RECT 551.995 -27.365 552.325 -27.035 ;
        RECT 550.635 -27.365 550.965 -27.035 ;
        RECT 549.275 -27.365 549.605 -27.035 ;
        RECT 547.915 -27.365 548.245 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.24 -35.52 554.36 -35.2 ;
        RECT 553.355 -35.525 553.685 -35.195 ;
        RECT 551.995 -35.525 552.325 -35.195 ;
        RECT 550.635 -35.525 550.965 -35.195 ;
        RECT 549.275 -35.525 549.605 -35.195 ;
        RECT 547.915 -35.525 548.245 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 547.24 -26 558.44 -25.68 ;
        RECT 556.075 -26.005 556.405 -25.675 ;
        RECT 551.995 -26.005 552.325 -25.675 ;
        RECT 550.635 -26.005 550.965 -25.675 ;
        RECT 549.275 -26.005 549.605 -25.675 ;
        RECT 547.915 -26.005 548.245 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -30.08 568.64 -29.76 ;
        RECT 566.955 -30.085 567.285 -29.755 ;
        RECT 565.595 -30.085 565.925 -29.755 ;
        RECT 564.235 -30.085 564.565 -29.755 ;
        RECT 562.875 -30.085 563.205 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.12 -23.28 569.32 -22.96 ;
        RECT 566.955 -23.285 567.285 -22.955 ;
        RECT 565.595 -23.285 565.925 -22.955 ;
        RECT 564.235 -23.285 564.565 -22.955 ;
        RECT 562.875 -23.285 563.205 -22.955 ;
        RECT 558.795 -23.285 559.125 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 558.8 -27.36 569.32 -27.04 ;
        RECT 566.955 -27.365 567.285 -27.035 ;
        RECT 565.595 -27.365 565.925 -27.035 ;
        RECT 564.235 -27.365 564.565 -27.035 ;
        RECT 562.875 -27.365 563.205 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -35.52 569.32 -35.2 ;
        RECT 568.315 -35.525 568.645 -35.195 ;
        RECT 566.955 -35.525 567.285 -35.195 ;
        RECT 565.595 -35.525 565.925 -35.195 ;
        RECT 564.235 -35.525 564.565 -35.195 ;
        RECT 562.875 -35.525 563.205 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 562.2 -26 572.72 -25.68 ;
        RECT 571.035 -26.005 571.365 -25.675 ;
        RECT 566.955 -26.005 567.285 -25.675 ;
        RECT 565.595 -26.005 565.925 -25.675 ;
        RECT 564.235 -26.005 564.565 -25.675 ;
        RECT 562.875 -26.005 563.205 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.16 -30.08 583.6 -29.76 ;
        RECT 581.915 -30.085 582.245 -29.755 ;
        RECT 580.555 -30.085 580.885 -29.755 ;
        RECT 579.195 -30.085 579.525 -29.755 ;
        RECT 577.835 -30.085 578.165 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.08 -23.28 584.28 -22.96 ;
        RECT 581.915 -23.285 582.245 -22.955 ;
        RECT 580.555 -23.285 580.885 -22.955 ;
        RECT 579.195 -23.285 579.525 -22.955 ;
        RECT 577.835 -23.285 578.165 -22.955 ;
        RECT 573.755 -23.285 574.085 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 573.76 -27.36 584.28 -27.04 ;
        RECT 581.915 -27.365 582.245 -27.035 ;
        RECT 580.555 -27.365 580.885 -27.035 ;
        RECT 579.195 -27.365 579.525 -27.035 ;
        RECT 577.835 -27.365 578.165 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.16 -35.52 584.28 -35.2 ;
        RECT 583.275 -35.525 583.605 -35.195 ;
        RECT 581.915 -35.525 582.245 -35.195 ;
        RECT 580.555 -35.525 580.885 -35.195 ;
        RECT 579.195 -35.525 579.525 -35.195 ;
        RECT 577.835 -35.525 578.165 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 577.16 -26 587.68 -25.68 ;
        RECT 585.995 -26.005 586.325 -25.675 ;
        RECT 581.915 -26.005 582.245 -25.675 ;
        RECT 580.555 -26.005 580.885 -25.675 ;
        RECT 579.195 -26.005 579.525 -25.675 ;
        RECT 577.835 -26.005 578.165 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.12 -30.08 598.56 -29.76 ;
        RECT 596.875 -30.085 597.205 -29.755 ;
        RECT 595.515 -30.085 595.845 -29.755 ;
        RECT 594.155 -30.085 594.485 -29.755 ;
        RECT 592.795 -30.085 593.125 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.04 -23.28 599.24 -22.96 ;
        RECT 596.875 -23.285 597.205 -22.955 ;
        RECT 595.515 -23.285 595.845 -22.955 ;
        RECT 594.155 -23.285 594.485 -22.955 ;
        RECT 592.795 -23.285 593.125 -22.955 ;
        RECT 588.715 -23.285 589.045 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 588.72 -27.36 599.24 -27.04 ;
        RECT 596.875 -27.365 597.205 -27.035 ;
        RECT 595.515 -27.365 595.845 -27.035 ;
        RECT 594.155 -27.365 594.485 -27.035 ;
        RECT 592.795 -27.365 593.125 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.12 -35.52 599.24 -35.2 ;
        RECT 598.235 -35.525 598.565 -35.195 ;
        RECT 596.875 -35.525 597.205 -35.195 ;
        RECT 595.515 -35.525 595.845 -35.195 ;
        RECT 594.155 -35.525 594.485 -35.195 ;
        RECT 592.795 -35.525 593.125 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 592.12 -26 602.64 -25.68 ;
        RECT 600.955 -26.005 601.285 -25.675 ;
        RECT 596.875 -26.005 597.205 -25.675 ;
        RECT 595.515 -26.005 595.845 -25.675 ;
        RECT 594.155 -26.005 594.485 -25.675 ;
        RECT 592.795 -26.005 593.125 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.08 -30.08 613.52 -29.76 ;
        RECT 611.835 -30.085 612.165 -29.755 ;
        RECT 610.475 -30.085 610.805 -29.755 ;
        RECT 609.115 -30.085 609.445 -29.755 ;
        RECT 607.755 -30.085 608.085 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 602.32 -23.28 614.2 -22.96 ;
        RECT 611.835 -23.285 612.165 -22.955 ;
        RECT 610.475 -23.285 610.805 -22.955 ;
        RECT 609.115 -23.285 609.445 -22.955 ;
        RECT 607.755 -23.285 608.085 -22.955 ;
        RECT 603.675 -23.285 604.005 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 603 -27.36 614.2 -27.04 ;
        RECT 611.835 -27.365 612.165 -27.035 ;
        RECT 610.475 -27.365 610.805 -27.035 ;
        RECT 609.115 -27.365 609.445 -27.035 ;
        RECT 607.755 -27.365 608.085 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.08 -35.52 614.2 -35.2 ;
        RECT 613.195 -35.525 613.525 -35.195 ;
        RECT 611.835 -35.525 612.165 -35.195 ;
        RECT 610.475 -35.525 610.805 -35.195 ;
        RECT 609.115 -35.525 609.445 -35.195 ;
        RECT 607.755 -35.525 608.085 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 607.08 -26 617.6 -25.68 ;
        RECT 615.915 -26.005 616.245 -25.675 ;
        RECT 611.835 -26.005 612.165 -25.675 ;
        RECT 610.475 -26.005 610.805 -25.675 ;
        RECT 609.115 -26.005 609.445 -25.675 ;
        RECT 607.755 -26.005 608.085 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.04 -30.08 628.48 -29.76 ;
        RECT 626.795 -30.085 627.125 -29.755 ;
        RECT 625.435 -30.085 625.765 -29.755 ;
        RECT 624.075 -30.085 624.405 -29.755 ;
        RECT 622.715 -30.085 623.045 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.28 -23.28 629.16 -22.96 ;
        RECT 626.795 -23.285 627.125 -22.955 ;
        RECT 625.435 -23.285 625.765 -22.955 ;
        RECT 624.075 -23.285 624.405 -22.955 ;
        RECT 622.715 -23.285 623.045 -22.955 ;
        RECT 618.635 -23.285 618.965 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 617.96 -27.36 629.16 -27.04 ;
        RECT 626.795 -27.365 627.125 -27.035 ;
        RECT 625.435 -27.365 625.765 -27.035 ;
        RECT 624.075 -27.365 624.405 -27.035 ;
        RECT 622.715 -27.365 623.045 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.04 -35.52 629.16 -35.2 ;
        RECT 628.155 -35.525 628.485 -35.195 ;
        RECT 626.795 -35.525 627.125 -35.195 ;
        RECT 625.435 -35.525 625.765 -35.195 ;
        RECT 624.075 -35.525 624.405 -35.195 ;
        RECT 622.715 -35.525 623.045 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 622.04 -26 632.56 -25.68 ;
        RECT 630.875 -26.005 631.205 -25.675 ;
        RECT 626.795 -26.005 627.125 -25.675 ;
        RECT 625.435 -26.005 625.765 -25.675 ;
        RECT 624.075 -26.005 624.405 -25.675 ;
        RECT 622.715 -26.005 623.045 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.24 -23.28 643.44 -22.96 ;
        RECT 641.755 -23.285 642.085 -22.955 ;
        RECT 640.395 -23.285 640.725 -22.955 ;
        RECT 639.035 -23.285 639.365 -22.955 ;
        RECT 637.675 -23.285 638.005 -22.955 ;
        RECT 633.595 -23.285 633.925 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 632.92 -27.36 643.44 -27.04 ;
        RECT 641.755 -27.365 642.085 -27.035 ;
        RECT 640.395 -27.365 640.725 -27.035 ;
        RECT 639.035 -27.365 639.365 -27.035 ;
        RECT 637.675 -27.365 638.005 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 637 -30.08 643.44 -29.76 ;
        RECT 641.755 -30.085 642.085 -29.755 ;
        RECT 640.395 -30.085 640.725 -29.755 ;
        RECT 639.035 -30.085 639.365 -29.755 ;
        RECT 637.675 -30.085 638.005 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 643.115 -35.525 643.445 -35.195 ;
        RECT 637 -35.52 643.445 -35.2 ;
        RECT 641.755 -35.525 642.085 -35.195 ;
        RECT 640.395 -35.525 640.725 -35.195 ;
        RECT 639.035 -35.525 639.365 -35.195 ;
        RECT 637.675 -35.525 638.005 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 637 -26 647.52 -25.68 ;
        RECT 645.835 -26.005 646.165 -25.675 ;
        RECT 641.755 -26.005 642.085 -25.675 ;
        RECT 640.395 -26.005 640.725 -25.675 ;
        RECT 639.035 -26.005 639.365 -25.675 ;
        RECT 637.675 -26.005 638.005 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.96 -30.08 657.72 -29.76 ;
        RECT 656.715 -30.085 657.045 -29.755 ;
        RECT 655.355 -30.085 655.685 -29.755 ;
        RECT 653.995 -30.085 654.325 -29.755 ;
        RECT 652.635 -30.085 652.965 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.2 -23.28 658.4 -22.96 ;
        RECT 656.715 -23.285 657.045 -22.955 ;
        RECT 655.355 -23.285 655.685 -22.955 ;
        RECT 653.995 -23.285 654.325 -22.955 ;
        RECT 652.635 -23.285 652.965 -22.955 ;
        RECT 648.555 -23.285 648.885 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 647.88 -27.36 658.4 -27.04 ;
        RECT 656.715 -27.365 657.045 -27.035 ;
        RECT 655.355 -27.365 655.685 -27.035 ;
        RECT 653.995 -27.365 654.325 -27.035 ;
        RECT 652.635 -27.365 652.965 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 658.075 -35.525 658.405 -35.195 ;
        RECT 651.96 -35.52 658.405 -35.2 ;
        RECT 656.715 -35.525 657.045 -35.195 ;
        RECT 655.355 -35.525 655.685 -35.195 ;
        RECT 653.995 -35.525 654.325 -35.195 ;
        RECT 652.635 -35.525 652.965 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 651.96 -26 662.48 -25.68 ;
        RECT 660.795 -26.005 661.125 -25.675 ;
        RECT 659.435 -26.005 659.765 -25.675 ;
        RECT 656.715 -26.005 657.045 -25.675 ;
        RECT 655.355 -26.005 655.685 -25.675 ;
        RECT 653.995 -26.005 654.325 -25.675 ;
        RECT 652.635 -26.005 652.965 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 666.92 -30.08 672.68 -29.76 ;
        RECT 671.675 -30.085 672.005 -29.755 ;
        RECT 670.315 -30.085 670.645 -29.755 ;
        RECT 668.955 -30.085 669.285 -29.755 ;
        RECT 667.595 -30.085 667.925 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.16 -23.28 673.36 -22.96 ;
        RECT 671.675 -23.285 672.005 -22.955 ;
        RECT 670.315 -23.285 670.645 -22.955 ;
        RECT 668.955 -23.285 669.285 -22.955 ;
        RECT 667.595 -23.285 667.925 -22.955 ;
        RECT 663.515 -23.285 663.845 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 662.84 -27.36 673.36 -27.04 ;
        RECT 671.675 -27.365 672.005 -27.035 ;
        RECT 670.315 -27.365 670.645 -27.035 ;
        RECT 668.955 -27.365 669.285 -27.035 ;
        RECT 667.595 -27.365 667.925 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 667.595 -35.525 667.925 -35.195 ;
        RECT 673.035 -35.525 673.365 -35.195 ;
        RECT 666.92 -35.52 673.365 -35.2 ;
        RECT 671.675 -35.525 672.005 -35.195 ;
        RECT 670.315 -35.525 670.645 -35.195 ;
        RECT 668.955 -35.525 669.285 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -23.28 2.88 -22.96 ;
        RECT 1.195 -23.285 1.525 -22.955 ;
        RECT -0.165 -23.285 0.165 -22.955 ;
        RECT -1.525 -23.285 -1.195 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -35.525 5.605 -35.195 ;
        RECT -1.525 -35.52 5.605 -35.2 ;
        RECT 3.915 -35.525 4.245 -35.195 ;
        RECT 2.555 -35.525 2.885 -35.195 ;
        RECT 1.195 -35.525 1.525 -35.195 ;
        RECT -0.165 -35.525 0.165 -35.195 ;
        RECT -1.525 -35.525 -1.195 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -30.08 17.16 -29.76 ;
        RECT 16.155 -30.085 16.485 -29.755 ;
        RECT 14.795 -30.085 15.125 -29.755 ;
        RECT 13.435 -30.085 13.765 -29.755 ;
        RECT 12.075 -30.085 12.405 -29.755 ;
        RECT 10.715 -30.085 11.045 -29.755 ;
        RECT 7.995 -30.085 8.325 -29.755 ;
        RECT 6.635 -30.085 6.965 -29.755 ;
        RECT 5.275 -30.085 5.605 -29.755 ;
        RECT 3.915 -30.085 4.245 -29.755 ;
        RECT 2.555 -30.085 2.885 -29.755 ;
        RECT 1.195 -30.085 1.525 -29.755 ;
        RECT -0.165 -30.085 0.165 -29.755 ;
        RECT -1.525 -30.085 -1.195 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -23.28 17.84 -22.96 ;
        RECT 16.155 -23.285 16.485 -22.955 ;
        RECT 14.795 -23.285 15.125 -22.955 ;
        RECT 13.435 -23.285 13.765 -22.955 ;
        RECT 12.075 -23.285 12.405 -22.955 ;
        RECT 10.715 -23.285 11.045 -22.955 ;
        RECT 7.995 -23.285 8.325 -22.955 ;
        RECT 6.635 -23.285 6.965 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -27.36 17.84 -27.04 ;
        RECT 16.155 -27.365 16.485 -27.035 ;
        RECT 14.795 -27.365 15.125 -27.035 ;
        RECT 13.435 -27.365 13.765 -27.035 ;
        RECT 12.075 -27.365 12.405 -27.035 ;
        RECT 10.715 -27.365 11.045 -27.035 ;
        RECT 7.995 -27.365 8.325 -27.035 ;
        RECT 6.635 -27.365 6.965 -27.035 ;
        RECT 5.275 -27.365 5.605 -27.035 ;
        RECT 3.915 -27.365 4.245 -27.035 ;
        RECT 2.555 -27.365 2.885 -27.035 ;
        RECT 1.195 -27.365 1.525 -27.035 ;
        RECT -0.165 -27.365 0.165 -27.035 ;
        RECT -1.525 -27.365 -1.195 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -35.525 17.845 -35.195 ;
        RECT 10.715 -35.52 17.845 -35.2 ;
        RECT 16.155 -35.525 16.485 -35.195 ;
        RECT 14.795 -35.525 15.125 -35.195 ;
        RECT 13.435 -35.525 13.765 -35.195 ;
        RECT 12.075 -35.525 12.405 -35.195 ;
        RECT 10.715 -35.525 11.045 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 -26 21.92 -25.68 ;
        RECT 20.235 -26.005 20.565 -25.675 ;
        RECT 18.875 -26.005 19.205 -25.675 ;
        RECT 16.155 -26.005 16.485 -25.675 ;
        RECT 14.795 -26.005 15.125 -25.675 ;
        RECT 13.435 -26.005 13.765 -25.675 ;
        RECT 12.075 -26.005 12.405 -25.675 ;
        RECT 10.715 -26.005 11.045 -25.675 ;
        RECT 7.995 -26.005 8.325 -25.675 ;
        RECT 6.635 -26.005 6.965 -25.675 ;
        RECT 5.275 -26.005 5.605 -25.675 ;
        RECT 3.915 -26.005 4.245 -25.675 ;
        RECT 2.555 -26.005 2.885 -25.675 ;
        RECT 1.195 -26.005 1.525 -25.675 ;
        RECT -0.165 -26.005 0.165 -25.675 ;
        RECT -1.525 -26.005 -1.195 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.68 -30.08 32.12 -29.76 ;
        RECT 31.115 -30.085 31.445 -29.755 ;
        RECT 29.755 -30.085 30.085 -29.755 ;
        RECT 28.395 -30.085 28.725 -29.755 ;
        RECT 27.035 -30.085 27.365 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.6 -23.28 32.8 -22.96 ;
        RECT 31.115 -23.285 31.445 -22.955 ;
        RECT 29.755 -23.285 30.085 -22.955 ;
        RECT 28.395 -23.285 28.725 -22.955 ;
        RECT 27.035 -23.285 27.365 -22.955 ;
        RECT 25.675 -23.285 26.005 -22.955 ;
        RECT 22.955 -23.285 23.285 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.28 -27.36 32.8 -27.04 ;
        RECT 31.115 -27.365 31.445 -27.035 ;
        RECT 29.755 -27.365 30.085 -27.035 ;
        RECT 28.395 -27.365 28.725 -27.035 ;
        RECT 27.035 -27.365 27.365 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -35.525 32.805 -35.195 ;
        RECT 25.68 -35.52 32.805 -35.2 ;
        RECT 31.115 -35.525 31.445 -35.195 ;
        RECT 29.755 -35.525 30.085 -35.195 ;
        RECT 28.395 -35.525 28.725 -35.195 ;
        RECT 27.035 -35.525 27.365 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.68 -26 36.88 -25.68 ;
        RECT 35.195 -26.005 35.525 -25.675 ;
        RECT 33.835 -26.005 34.165 -25.675 ;
        RECT 31.115 -26.005 31.445 -25.675 ;
        RECT 29.755 -26.005 30.085 -25.675 ;
        RECT 28.395 -26.005 28.725 -25.675 ;
        RECT 27.035 -26.005 27.365 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.64 -30.08 47.08 -29.76 ;
        RECT 46.075 -30.085 46.405 -29.755 ;
        RECT 44.715 -30.085 45.045 -29.755 ;
        RECT 43.355 -30.085 43.685 -29.755 ;
        RECT 41.995 -30.085 42.325 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.56 -23.28 47.76 -22.96 ;
        RECT 46.075 -23.285 46.405 -22.955 ;
        RECT 44.715 -23.285 45.045 -22.955 ;
        RECT 43.355 -23.285 43.685 -22.955 ;
        RECT 41.995 -23.285 42.325 -22.955 ;
        RECT 40.635 -23.285 40.965 -22.955 ;
        RECT 37.915 -23.285 38.245 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.24 -27.36 47.76 -27.04 ;
        RECT 46.075 -27.365 46.405 -27.035 ;
        RECT 44.715 -27.365 45.045 -27.035 ;
        RECT 43.355 -27.365 43.685 -27.035 ;
        RECT 41.995 -27.365 42.325 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 -35.525 47.765 -35.195 ;
        RECT 40.64 -35.52 47.765 -35.2 ;
        RECT 46.075 -35.525 46.405 -35.195 ;
        RECT 44.715 -35.525 45.045 -35.195 ;
        RECT 43.355 -35.525 43.685 -35.195 ;
        RECT 41.995 -35.525 42.325 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.64 -26 51.84 -25.68 ;
        RECT 50.155 -26.005 50.485 -25.675 ;
        RECT 48.795 -26.005 49.125 -25.675 ;
        RECT 46.075 -26.005 46.405 -25.675 ;
        RECT 44.715 -26.005 45.045 -25.675 ;
        RECT 43.355 -26.005 43.685 -25.675 ;
        RECT 41.995 -26.005 42.325 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.6 -30.08 62.04 -29.76 ;
        RECT 61.035 -30.085 61.365 -29.755 ;
        RECT 59.675 -30.085 60.005 -29.755 ;
        RECT 58.315 -30.085 58.645 -29.755 ;
        RECT 56.955 -30.085 57.285 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.52 -23.28 62.72 -22.96 ;
        RECT 61.035 -23.285 61.365 -22.955 ;
        RECT 59.675 -23.285 60.005 -22.955 ;
        RECT 58.315 -23.285 58.645 -22.955 ;
        RECT 56.955 -23.285 57.285 -22.955 ;
        RECT 55.595 -23.285 55.925 -22.955 ;
        RECT 52.875 -23.285 53.205 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.2 -27.36 62.72 -27.04 ;
        RECT 61.035 -27.365 61.365 -27.035 ;
        RECT 59.675 -27.365 60.005 -27.035 ;
        RECT 58.315 -27.365 58.645 -27.035 ;
        RECT 56.955 -27.365 57.285 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -35.525 62.725 -35.195 ;
        RECT 55.6 -35.52 62.725 -35.2 ;
        RECT 61.035 -35.525 61.365 -35.195 ;
        RECT 59.675 -35.525 60.005 -35.195 ;
        RECT 58.315 -35.525 58.645 -35.195 ;
        RECT 56.955 -35.525 57.285 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.6 -26 66.12 -25.68 ;
        RECT 65.115 -26.005 65.445 -25.675 ;
        RECT 63.755 -26.005 64.085 -25.675 ;
        RECT 61.035 -26.005 61.365 -25.675 ;
        RECT 59.675 -26.005 60.005 -25.675 ;
        RECT 58.315 -26.005 58.645 -25.675 ;
        RECT 56.955 -26.005 57.285 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.56 -30.08 77 -29.76 ;
        RECT 75.995 -30.085 76.325 -29.755 ;
        RECT 74.635 -30.085 74.965 -29.755 ;
        RECT 73.275 -30.085 73.605 -29.755 ;
        RECT 71.915 -30.085 72.245 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.48 -23.28 77.68 -22.96 ;
        RECT 75.995 -23.285 76.325 -22.955 ;
        RECT 74.635 -23.285 74.965 -22.955 ;
        RECT 73.275 -23.285 73.605 -22.955 ;
        RECT 71.915 -23.285 72.245 -22.955 ;
        RECT 70.555 -23.285 70.885 -22.955 ;
        RECT 67.835 -23.285 68.165 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.16 -27.36 77.68 -27.04 ;
        RECT 75.995 -27.365 76.325 -27.035 ;
        RECT 74.635 -27.365 74.965 -27.035 ;
        RECT 73.275 -27.365 73.605 -27.035 ;
        RECT 71.915 -27.365 72.245 -27.035 ;
        RECT 67.835 -27.365 68.165 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -35.525 77.685 -35.195 ;
        RECT 70.56 -35.52 77.685 -35.2 ;
        RECT 75.995 -35.525 76.325 -35.195 ;
        RECT 74.635 -35.525 74.965 -35.195 ;
        RECT 73.275 -35.525 73.605 -35.195 ;
        RECT 71.915 -35.525 72.245 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.56 -26 81.08 -25.68 ;
        RECT 80.075 -26.005 80.405 -25.675 ;
        RECT 78.715 -26.005 79.045 -25.675 ;
        RECT 75.995 -26.005 76.325 -25.675 ;
        RECT 74.635 -26.005 74.965 -25.675 ;
        RECT 73.275 -26.005 73.605 -25.675 ;
        RECT 71.915 -26.005 72.245 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.52 -30.08 91.96 -29.76 ;
        RECT 90.955 -30.085 91.285 -29.755 ;
        RECT 89.595 -30.085 89.925 -29.755 ;
        RECT 88.235 -30.085 88.565 -29.755 ;
        RECT 86.875 -30.085 87.205 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 -23.28 92.64 -22.96 ;
        RECT 90.955 -23.285 91.285 -22.955 ;
        RECT 89.595 -23.285 89.925 -22.955 ;
        RECT 88.235 -23.285 88.565 -22.955 ;
        RECT 86.875 -23.285 87.205 -22.955 ;
        RECT 85.515 -23.285 85.845 -22.955 ;
        RECT 82.795 -23.285 83.125 -22.955 ;
        RECT 81.435 -23.285 81.765 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.12 -27.36 92.64 -27.04 ;
        RECT 90.955 -27.365 91.285 -27.035 ;
        RECT 89.595 -27.365 89.925 -27.035 ;
        RECT 88.235 -27.365 88.565 -27.035 ;
        RECT 86.875 -27.365 87.205 -27.035 ;
        RECT 82.795 -27.365 83.125 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -35.525 92.645 -35.195 ;
        RECT 85.52 -35.52 92.645 -35.2 ;
        RECT 90.955 -35.525 91.285 -35.195 ;
        RECT 89.595 -35.525 89.925 -35.195 ;
        RECT 88.235 -35.525 88.565 -35.195 ;
        RECT 86.875 -35.525 87.205 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.52 -26 96.04 -25.68 ;
        RECT 93.675 -26.005 94.005 -25.675 ;
        RECT 90.955 -26.005 91.285 -25.675 ;
        RECT 89.595 -26.005 89.925 -25.675 ;
        RECT 88.235 -26.005 88.565 -25.675 ;
        RECT 86.875 -26.005 87.205 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.48 -30.08 106.92 -29.76 ;
        RECT 105.915 -30.085 106.245 -29.755 ;
        RECT 104.555 -30.085 104.885 -29.755 ;
        RECT 103.195 -30.085 103.525 -29.755 ;
        RECT 101.835 -30.085 102.165 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.72 -23.28 107.6 -22.96 ;
        RECT 105.915 -23.285 106.245 -22.955 ;
        RECT 104.555 -23.285 104.885 -22.955 ;
        RECT 103.195 -23.285 103.525 -22.955 ;
        RECT 101.835 -23.285 102.165 -22.955 ;
        RECT 100.475 -23.285 100.805 -22.955 ;
        RECT 97.755 -23.285 98.085 -22.955 ;
        RECT 96.395 -23.285 96.725 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.4 -27.36 107.6 -27.04 ;
        RECT 105.915 -27.365 106.245 -27.035 ;
        RECT 104.555 -27.365 104.885 -27.035 ;
        RECT 103.195 -27.365 103.525 -27.035 ;
        RECT 101.835 -27.365 102.165 -27.035 ;
        RECT 97.755 -27.365 98.085 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 -35.525 107.605 -35.195 ;
        RECT 100.48 -35.52 107.605 -35.2 ;
        RECT 105.915 -35.525 106.245 -35.195 ;
        RECT 104.555 -35.525 104.885 -35.195 ;
        RECT 103.195 -35.525 103.525 -35.195 ;
        RECT 101.835 -35.525 102.165 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.48 -26 111 -25.68 ;
        RECT 108.635 -26.005 108.965 -25.675 ;
        RECT 105.915 -26.005 106.245 -25.675 ;
        RECT 104.555 -26.005 104.885 -25.675 ;
        RECT 103.195 -26.005 103.525 -25.675 ;
        RECT 101.835 -26.005 102.165 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.44 -30.08 121.88 -29.76 ;
        RECT 120.875 -30.085 121.205 -29.755 ;
        RECT 119.515 -30.085 119.845 -29.755 ;
        RECT 118.155 -30.085 118.485 -29.755 ;
        RECT 116.795 -30.085 117.125 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.68 -23.28 122.56 -22.96 ;
        RECT 120.875 -23.285 121.205 -22.955 ;
        RECT 119.515 -23.285 119.845 -22.955 ;
        RECT 118.155 -23.285 118.485 -22.955 ;
        RECT 116.795 -23.285 117.125 -22.955 ;
        RECT 115.435 -23.285 115.765 -22.955 ;
        RECT 112.715 -23.285 113.045 -22.955 ;
        RECT 111.355 -23.285 111.685 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.36 -27.36 122.56 -27.04 ;
        RECT 120.875 -27.365 121.205 -27.035 ;
        RECT 119.515 -27.365 119.845 -27.035 ;
        RECT 118.155 -27.365 118.485 -27.035 ;
        RECT 116.795 -27.365 117.125 -27.035 ;
        RECT 112.715 -27.365 113.045 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 -35.525 122.565 -35.195 ;
        RECT 115.44 -35.52 122.565 -35.2 ;
        RECT 120.875 -35.525 121.205 -35.195 ;
        RECT 119.515 -35.525 119.845 -35.195 ;
        RECT 118.155 -35.525 118.485 -35.195 ;
        RECT 116.795 -35.525 117.125 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.44 -26 125.96 -25.68 ;
        RECT 123.595 -26.005 123.925 -25.675 ;
        RECT 120.875 -26.005 121.205 -25.675 ;
        RECT 119.515 -26.005 119.845 -25.675 ;
        RECT 118.155 -26.005 118.485 -25.675 ;
        RECT 116.795 -26.005 117.125 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.64 -23.28 136.84 -22.96 ;
        RECT 134.475 -23.285 134.805 -22.955 ;
        RECT 133.115 -23.285 133.445 -22.955 ;
        RECT 131.755 -23.285 132.085 -22.955 ;
        RECT 130.395 -23.285 130.725 -22.955 ;
        RECT 127.675 -23.285 128.005 -22.955 ;
        RECT 126.315 -23.285 126.645 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.32 -27.36 136.84 -27.04 ;
        RECT 134.475 -27.365 134.805 -27.035 ;
        RECT 133.115 -27.365 133.445 -27.035 ;
        RECT 131.755 -27.365 132.085 -27.035 ;
        RECT 127.675 -27.365 128.005 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.4 -30.08 136.84 -29.76 ;
        RECT 134.475 -30.085 134.805 -29.755 ;
        RECT 133.115 -30.085 133.445 -29.755 ;
        RECT 131.755 -30.085 132.085 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.4 -35.52 136.84 -35.2 ;
        RECT 135.835 -35.525 136.165 -35.195 ;
        RECT 134.475 -35.525 134.805 -35.195 ;
        RECT 133.115 -35.525 133.445 -35.195 ;
        RECT 131.755 -35.525 132.085 -35.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.4 -26 140.92 -25.68 ;
        RECT 138.555 -26.005 138.885 -25.675 ;
        RECT 134.475 -26.005 134.805 -25.675 ;
        RECT 133.115 -26.005 133.445 -25.675 ;
        RECT 131.755 -26.005 132.085 -25.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.36 -30.08 151.12 -29.76 ;
        RECT 149.435 -30.085 149.765 -29.755 ;
        RECT 148.075 -30.085 148.405 -29.755 ;
        RECT 146.715 -30.085 147.045 -29.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -23.28 151.8 -22.96 ;
        RECT 149.435 -23.285 149.765 -22.955 ;
        RECT 148.075 -23.285 148.405 -22.955 ;
        RECT 146.715 -23.285 147.045 -22.955 ;
        RECT 145.355 -23.285 145.685 -22.955 ;
        RECT 142.635 -23.285 142.965 -22.955 ;
        RECT 141.275 -23.285 141.605 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -27.365 148.405 -27.035 ;
        RECT 146.715 -27.365 147.045 -27.035 ;
        RECT 142.635 -27.365 142.965 -27.035 ;
        RECT 141.28 -27.36 151.8 -27.04 ;
        RECT 149.435 -27.365 149.765 -27.035 ;
    END
  END vss
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.26 -35.475 6.58 -35.145 ;
        RECT 6.28 -35.495 6.56 -35.125 ;
    END
  END dout[0]
  PIN dout[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.76 -35.47 379.08 -35.15 ;
    END
  END dout[100]
  PIN dout[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.02 -35.47 380.34 -35.15 ;
    END
  END dout[101]
  PIN dout[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.14 -35.475 391.46 -35.145 ;
        RECT 391.16 -35.495 391.44 -35.125 ;
    END
  END dout[102]
  PIN dout[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.4 -35.47 392.72 -35.15 ;
    END
  END dout[103]
  PIN dout[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.66 -35.47 393.98 -35.15 ;
    END
  END dout[104]
  PIN dout[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.92 -35.47 395.24 -35.15 ;
    END
  END dout[105]
  PIN dout[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.04 -35.475 406.36 -35.145 ;
        RECT 406.06 -35.495 406.34 -35.125 ;
    END
  END dout[106]
  PIN dout[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.3 -35.47 407.62 -35.15 ;
    END
  END dout[107]
  PIN dout[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.56 -35.47 408.88 -35.15 ;
    END
  END dout[108]
  PIN dout[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.82 -35.47 410.14 -35.15 ;
    END
  END dout[109]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.44 -35.475 48.76 -35.145 ;
        RECT 48.46 -35.495 48.74 -35.125 ;
    END
  END dout[10]
  PIN dout[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.94 -35.475 421.26 -35.145 ;
        RECT 420.96 -35.495 421.24 -35.125 ;
    END
  END dout[110]
  PIN dout[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.2 -35.47 422.52 -35.15 ;
    END
  END dout[111]
  PIN dout[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.46 -35.47 423.78 -35.15 ;
    END
  END dout[112]
  PIN dout[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.72 -35.47 425.04 -35.15 ;
    END
  END dout[113]
  PIN dout[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.84 -35.475 436.16 -35.145 ;
        RECT 435.86 -35.495 436.14 -35.125 ;
    END
  END dout[114]
  PIN dout[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.1 -35.47 437.42 -35.15 ;
    END
  END dout[115]
  PIN dout[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.36 -35.47 438.68 -35.15 ;
    END
  END dout[116]
  PIN dout[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.62 -35.47 439.94 -35.15 ;
    END
  END dout[117]
  PIN dout[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.74 -35.475 451.06 -35.145 ;
        RECT 450.76 -35.495 451.04 -35.125 ;
    END
  END dout[118]
  PIN dout[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452 -35.47 452.32 -35.15 ;
    END
  END dout[119]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.7 -35.47 50.02 -35.15 ;
    END
  END dout[11]
  PIN dout[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.26 -35.47 453.58 -35.15 ;
    END
  END dout[120]
  PIN dout[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.52 -35.47 454.84 -35.15 ;
    END
  END dout[121]
  PIN dout[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.64 -35.475 465.96 -35.145 ;
        RECT 465.66 -35.495 465.94 -35.125 ;
    END
  END dout[122]
  PIN dout[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.9 -35.47 467.22 -35.15 ;
    END
  END dout[123]
  PIN dout[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.16 -35.47 468.48 -35.15 ;
    END
  END dout[124]
  PIN dout[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.42 -35.47 469.74 -35.15 ;
    END
  END dout[125]
  PIN dout[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.54 -35.475 480.86 -35.145 ;
        RECT 480.56 -35.495 480.84 -35.125 ;
    END
  END dout[126]
  PIN dout[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.8 -35.47 482.12 -35.15 ;
    END
  END dout[127]
  PIN dout[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.06 -35.47 483.38 -35.15 ;
    END
  END dout[128]
  PIN dout[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.32 -35.47 484.64 -35.15 ;
    END
  END dout[129]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.96 -35.47 51.28 -35.15 ;
    END
  END dout[12]
  PIN dout[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.44 -35.475 495.76 -35.145 ;
        RECT 495.46 -35.495 495.74 -35.125 ;
    END
  END dout[130]
  PIN dout[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.7 -35.47 497.02 -35.15 ;
    END
  END dout[131]
  PIN dout[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.96 -35.47 498.28 -35.15 ;
    END
  END dout[132]
  PIN dout[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.22 -35.47 499.54 -35.15 ;
    END
  END dout[133]
  PIN dout[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.34 -35.475 510.66 -35.145 ;
        RECT 510.36 -35.495 510.64 -35.125 ;
    END
  END dout[134]
  PIN dout[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.6 -35.47 511.92 -35.15 ;
    END
  END dout[135]
  PIN dout[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.86 -35.47 513.18 -35.15 ;
    END
  END dout[136]
  PIN dout[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.12 -35.47 514.44 -35.15 ;
    END
  END dout[137]
  PIN dout[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.24 -35.475 525.56 -35.145 ;
        RECT 525.26 -35.495 525.54 -35.125 ;
    END
  END dout[138]
  PIN dout[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.5 -35.47 526.82 -35.15 ;
    END
  END dout[139]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.22 -35.47 52.54 -35.15 ;
    END
  END dout[13]
  PIN dout[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.76 -35.47 528.08 -35.15 ;
    END
  END dout[140]
  PIN dout[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.02 -35.47 529.34 -35.15 ;
    END
  END dout[141]
  PIN dout[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.14 -35.475 540.46 -35.145 ;
        RECT 540.16 -35.495 540.44 -35.125 ;
    END
  END dout[142]
  PIN dout[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.4 -35.47 541.72 -35.15 ;
    END
  END dout[143]
  PIN dout[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.66 -35.47 542.98 -35.15 ;
    END
  END dout[144]
  PIN dout[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.92 -35.47 544.24 -35.15 ;
    END
  END dout[145]
  PIN dout[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.04 -35.475 555.36 -35.145 ;
        RECT 555.06 -35.495 555.34 -35.125 ;
    END
  END dout[146]
  PIN dout[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.3 -35.47 556.62 -35.15 ;
    END
  END dout[147]
  PIN dout[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.56 -35.47 557.88 -35.15 ;
    END
  END dout[148]
  PIN dout[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.82 -35.47 559.14 -35.15 ;
    END
  END dout[149]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.34 -35.475 63.66 -35.145 ;
        RECT 63.36 -35.495 63.64 -35.125 ;
    END
  END dout[14]
  PIN dout[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.94 -35.475 570.26 -35.145 ;
        RECT 569.96 -35.495 570.24 -35.125 ;
    END
  END dout[150]
  PIN dout[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.2 -35.47 571.52 -35.15 ;
    END
  END dout[151]
  PIN dout[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.46 -35.47 572.78 -35.15 ;
    END
  END dout[152]
  PIN dout[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.72 -35.47 574.04 -35.15 ;
    END
  END dout[153]
  PIN dout[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.84 -35.475 585.16 -35.145 ;
        RECT 584.86 -35.495 585.14 -35.125 ;
    END
  END dout[154]
  PIN dout[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.1 -35.47 586.42 -35.15 ;
    END
  END dout[155]
  PIN dout[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.36 -35.47 587.68 -35.15 ;
    END
  END dout[156]
  PIN dout[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.62 -35.47 588.94 -35.15 ;
    END
  END dout[157]
  PIN dout[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.74 -35.475 600.06 -35.145 ;
        RECT 599.76 -35.495 600.04 -35.125 ;
    END
  END dout[158]
  PIN dout[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601 -35.47 601.32 -35.15 ;
    END
  END dout[159]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.6 -35.47 64.92 -35.15 ;
    END
  END dout[15]
  PIN dout[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.26 -35.47 602.58 -35.15 ;
    END
  END dout[160]
  PIN dout[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.52 -35.47 603.84 -35.15 ;
    END
  END dout[161]
  PIN dout[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.64 -35.475 614.96 -35.145 ;
        RECT 614.66 -35.495 614.94 -35.125 ;
    END
  END dout[162]
  PIN dout[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.9 -35.47 616.22 -35.15 ;
    END
  END dout[163]
  PIN dout[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.16 -35.47 617.48 -35.15 ;
    END
  END dout[164]
  PIN dout[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.42 -35.47 618.74 -35.15 ;
    END
  END dout[165]
  PIN dout[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.54 -35.475 629.86 -35.145 ;
        RECT 629.56 -35.495 629.84 -35.125 ;
    END
  END dout[166]
  PIN dout[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.8 -35.47 631.12 -35.15 ;
    END
  END dout[167]
  PIN dout[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.06 -35.47 632.38 -35.15 ;
    END
  END dout[168]
  PIN dout[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.32 -35.47 633.64 -35.15 ;
    END
  END dout[169]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.86 -35.47 66.18 -35.15 ;
    END
  END dout[16]
  PIN dout[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.44 -35.475 644.76 -35.145 ;
        RECT 644.46 -35.495 644.74 -35.125 ;
    END
  END dout[170]
  PIN dout[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.7 -35.47 646.02 -35.15 ;
    END
  END dout[171]
  PIN dout[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.96 -35.47 647.28 -35.15 ;
    END
  END dout[172]
  PIN dout[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.22 -35.47 648.54 -35.15 ;
    END
  END dout[173]
  PIN dout[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.34 -35.475 659.66 -35.145 ;
        RECT 659.36 -35.495 659.64 -35.125 ;
    END
  END dout[174]
  PIN dout[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.6 -35.47 660.92 -35.15 ;
    END
  END dout[175]
  PIN dout[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.86 -35.47 662.18 -35.15 ;
    END
  END dout[176]
  PIN dout[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.12 -35.47 663.44 -35.15 ;
    END
  END dout[177]
  PIN dout[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.24 -35.475 674.56 -35.145 ;
        RECT 674.26 -35.495 674.54 -35.125 ;
    END
  END dout[178]
  PIN dout[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.5 -35.47 675.82 -35.15 ;
    END
  END dout[179]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.12 -35.47 67.44 -35.15 ;
    END
  END dout[17]
  PIN dout[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.76 -35.47 677.08 -35.15 ;
    END
  END dout[180]
  PIN dout[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.02 -35.47 678.34 -35.15 ;
    END
  END dout[181]
  PIN dout[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.14 -35.475 689.46 -35.145 ;
        RECT 689.16 -35.495 689.44 -35.125 ;
    END
  END dout[182]
  PIN dout[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.4 -35.47 690.72 -35.15 ;
    END
  END dout[183]
  PIN dout[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.66 -35.47 691.98 -35.15 ;
    END
  END dout[184]
  PIN dout[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.92 -35.47 693.24 -35.15 ;
    END
  END dout[185]
  PIN dout[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.04 -35.475 704.36 -35.145 ;
        RECT 704.06 -35.495 704.34 -35.125 ;
    END
  END dout[186]
  PIN dout[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.3 -35.47 705.62 -35.15 ;
    END
  END dout[187]
  PIN dout[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.56 -35.47 706.88 -35.15 ;
    END
  END dout[188]
  PIN dout[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.82 -35.47 708.14 -35.15 ;
    END
  END dout[189]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.24 -35.475 78.56 -35.145 ;
        RECT 78.26 -35.495 78.54 -35.125 ;
    END
  END dout[18]
  PIN dout[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.94 -35.475 719.26 -35.145 ;
        RECT 718.96 -35.495 719.24 -35.125 ;
    END
  END dout[190]
  PIN dout[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.2 -35.47 720.52 -35.15 ;
    END
  END dout[191]
  PIN dout[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.46 -35.47 721.78 -35.15 ;
    END
  END dout[192]
  PIN dout[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.72 -35.47 723.04 -35.15 ;
    END
  END dout[193]
  PIN dout[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.84 -35.475 734.16 -35.145 ;
        RECT 733.86 -35.495 734.14 -35.125 ;
    END
  END dout[194]
  PIN dout[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.1 -35.47 735.42 -35.15 ;
    END
  END dout[195]
  PIN dout[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.36 -35.47 736.68 -35.15 ;
    END
  END dout[196]
  PIN dout[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.62 -35.47 737.94 -35.15 ;
    END
  END dout[197]
  PIN dout[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.74 -35.475 749.06 -35.145 ;
        RECT 748.76 -35.495 749.04 -35.125 ;
    END
  END dout[198]
  PIN dout[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750 -35.47 750.32 -35.15 ;
    END
  END dout[199]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.5 -35.47 79.82 -35.15 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 -35.47 7.84 -35.15 ;
    END
  END dout[1]
  PIN dout[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.26 -35.47 751.58 -35.15 ;
    END
  END dout[200]
  PIN dout[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.52 -35.47 752.84 -35.15 ;
    END
  END dout[201]
  PIN dout[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.64 -35.475 763.96 -35.145 ;
        RECT 763.66 -35.495 763.94 -35.125 ;
    END
  END dout[202]
  PIN dout[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.9 -35.47 765.22 -35.15 ;
    END
  END dout[203]
  PIN dout[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.16 -35.47 766.48 -35.15 ;
    END
  END dout[204]
  PIN dout[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.42 -35.47 767.74 -35.15 ;
    END
  END dout[205]
  PIN dout[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.54 -35.475 778.86 -35.145 ;
        RECT 778.56 -35.495 778.84 -35.125 ;
    END
  END dout[206]
  PIN dout[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.8 -35.47 780.12 -35.15 ;
    END
  END dout[207]
  PIN dout[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.06 -35.47 781.38 -35.15 ;
    END
  END dout[208]
  PIN dout[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.32 -35.47 782.64 -35.15 ;
    END
  END dout[209]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.76 -35.47 81.08 -35.15 ;
    END
  END dout[20]
  PIN dout[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.44 -35.475 793.76 -35.145 ;
        RECT 793.46 -35.495 793.74 -35.125 ;
    END
  END dout[210]
  PIN dout[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.7 -35.47 795.02 -35.15 ;
    END
  END dout[211]
  PIN dout[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.96 -35.47 796.28 -35.15 ;
    END
  END dout[212]
  PIN dout[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.22 -35.47 797.54 -35.15 ;
    END
  END dout[213]
  PIN dout[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.34 -35.475 808.66 -35.145 ;
        RECT 808.36 -35.495 808.64 -35.125 ;
    END
  END dout[214]
  PIN dout[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.6 -35.47 809.92 -35.15 ;
    END
  END dout[215]
  PIN dout[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.86 -35.47 811.18 -35.15 ;
    END
  END dout[216]
  PIN dout[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.12 -35.47 812.44 -35.15 ;
    END
  END dout[217]
  PIN dout[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.24 -35.475 823.56 -35.145 ;
        RECT 823.26 -35.495 823.54 -35.125 ;
    END
  END dout[218]
  PIN dout[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.5 -35.47 824.82 -35.15 ;
    END
  END dout[219]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.02 -35.47 82.34 -35.15 ;
    END
  END dout[21]
  PIN dout[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.76 -35.47 826.08 -35.15 ;
    END
  END dout[220]
  PIN dout[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.02 -35.47 827.34 -35.15 ;
    END
  END dout[221]
  PIN dout[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.14 -35.475 838.46 -35.145 ;
        RECT 838.16 -35.495 838.44 -35.125 ;
    END
  END dout[222]
  PIN dout[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.4 -35.47 839.72 -35.15 ;
    END
  END dout[223]
  PIN dout[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.66 -35.47 840.98 -35.15 ;
    END
  END dout[224]
  PIN dout[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.92 -35.47 842.24 -35.15 ;
    END
  END dout[225]
  PIN dout[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.04 -35.475 853.36 -35.145 ;
        RECT 853.06 -35.495 853.34 -35.125 ;
    END
  END dout[226]
  PIN dout[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.3 -35.47 854.62 -35.15 ;
    END
  END dout[227]
  PIN dout[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.56 -35.47 855.88 -35.15 ;
    END
  END dout[228]
  PIN dout[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.82 -35.47 857.14 -35.15 ;
    END
  END dout[229]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.14 -35.475 93.46 -35.145 ;
        RECT 93.16 -35.495 93.44 -35.125 ;
    END
  END dout[22]
  PIN dout[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.94 -35.475 868.26 -35.145 ;
        RECT 867.96 -35.495 868.24 -35.125 ;
    END
  END dout[230]
  PIN dout[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.2 -35.47 869.52 -35.15 ;
    END
  END dout[231]
  PIN dout[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.46 -35.47 870.78 -35.15 ;
    END
  END dout[232]
  PIN dout[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.72 -35.47 872.04 -35.15 ;
    END
  END dout[233]
  PIN dout[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.84 -35.475 883.16 -35.145 ;
        RECT 882.86 -35.495 883.14 -35.125 ;
    END
  END dout[234]
  PIN dout[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.1 -35.47 884.42 -35.15 ;
    END
  END dout[235]
  PIN dout[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.36 -35.47 885.68 -35.15 ;
    END
  END dout[236]
  PIN dout[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.62 -35.47 886.94 -35.15 ;
    END
  END dout[237]
  PIN dout[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.74 -35.475 898.06 -35.145 ;
        RECT 897.76 -35.495 898.04 -35.125 ;
    END
  END dout[238]
  PIN dout[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899 -35.47 899.32 -35.15 ;
    END
  END dout[239]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.4 -35.47 94.72 -35.15 ;
    END
  END dout[23]
  PIN dout[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.26 -35.47 900.58 -35.15 ;
    END
  END dout[240]
  PIN dout[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.52 -35.47 901.84 -35.15 ;
    END
  END dout[241]
  PIN dout[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.64 -35.475 912.96 -35.145 ;
        RECT 912.66 -35.495 912.94 -35.125 ;
    END
  END dout[242]
  PIN dout[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.9 -35.47 914.22 -35.15 ;
    END
  END dout[243]
  PIN dout[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.16 -35.47 915.48 -35.15 ;
    END
  END dout[244]
  PIN dout[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.42 -35.47 916.74 -35.15 ;
    END
  END dout[245]
  PIN dout[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.54 -35.475 927.86 -35.145 ;
        RECT 927.56 -35.495 927.84 -35.125 ;
    END
  END dout[246]
  PIN dout[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.8 -35.47 929.12 -35.15 ;
    END
  END dout[247]
  PIN dout[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.06 -35.47 930.38 -35.15 ;
    END
  END dout[248]
  PIN dout[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.32 -35.47 931.64 -35.15 ;
    END
  END dout[249]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.66 -35.47 95.98 -35.15 ;
    END
  END dout[24]
  PIN dout[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.96 -35.475 945.28 -35.145 ;
        RECT 944.98 -35.495 945.26 -35.125 ;
    END
  END dout[250]
  PIN dout[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.22 -35.47 946.54 -35.15 ;
    END
  END dout[251]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.92 -35.47 97.24 -35.15 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.04 -35.475 108.36 -35.145 ;
        RECT 108.06 -35.495 108.34 -35.125 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.3 -35.47 109.62 -35.15 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.56 -35.47 110.88 -35.15 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.82 -35.47 112.14 -35.15 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.64 -35.475 18.96 -35.145 ;
        RECT 18.66 -35.495 18.94 -35.125 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.94 -35.475 123.26 -35.145 ;
        RECT 122.96 -35.495 123.24 -35.125 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.2 -35.47 124.52 -35.15 ;
    END
  END dout[31]
  PIN dout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.46 -35.47 125.78 -35.15 ;
    END
  END dout[32]
  PIN dout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.72 -35.47 127.04 -35.15 ;
    END
  END dout[33]
  PIN dout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.84 -35.475 138.16 -35.145 ;
        RECT 137.86 -35.495 138.14 -35.125 ;
    END
  END dout[34]
  PIN dout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.1 -35.47 139.42 -35.15 ;
    END
  END dout[35]
  PIN dout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.36 -35.47 140.68 -35.15 ;
    END
  END dout[36]
  PIN dout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.62 -35.47 141.94 -35.15 ;
    END
  END dout[37]
  PIN dout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.74 -35.475 153.06 -35.145 ;
        RECT 152.76 -35.495 153.04 -35.125 ;
    END
  END dout[38]
  PIN dout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154 -35.47 154.32 -35.15 ;
    END
  END dout[39]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.9 -35.47 20.22 -35.15 ;
    END
  END dout[3]
  PIN dout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.26 -35.47 155.58 -35.15 ;
    END
  END dout[40]
  PIN dout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.52 -35.47 156.84 -35.15 ;
    END
  END dout[41]
  PIN dout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.64 -35.475 167.96 -35.145 ;
        RECT 167.66 -35.495 167.94 -35.125 ;
    END
  END dout[42]
  PIN dout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.9 -35.47 169.22 -35.15 ;
    END
  END dout[43]
  PIN dout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.16 -35.47 170.48 -35.15 ;
    END
  END dout[44]
  PIN dout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.42 -35.47 171.74 -35.15 ;
    END
  END dout[45]
  PIN dout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.54 -35.475 182.86 -35.145 ;
        RECT 182.56 -35.495 182.84 -35.125 ;
    END
  END dout[46]
  PIN dout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.8 -35.47 184.12 -35.15 ;
    END
  END dout[47]
  PIN dout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.06 -35.47 185.38 -35.15 ;
    END
  END dout[48]
  PIN dout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.32 -35.47 186.64 -35.15 ;
    END
  END dout[49]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.16 -35.47 21.48 -35.15 ;
    END
  END dout[4]
  PIN dout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.44 -35.475 197.76 -35.145 ;
        RECT 197.46 -35.495 197.74 -35.125 ;
    END
  END dout[50]
  PIN dout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.7 -35.47 199.02 -35.15 ;
    END
  END dout[51]
  PIN dout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.96 -35.47 200.28 -35.15 ;
    END
  END dout[52]
  PIN dout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.22 -35.47 201.54 -35.15 ;
    END
  END dout[53]
  PIN dout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.34 -35.475 212.66 -35.145 ;
        RECT 212.36 -35.495 212.64 -35.125 ;
    END
  END dout[54]
  PIN dout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.6 -35.47 213.92 -35.15 ;
    END
  END dout[55]
  PIN dout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.86 -35.47 215.18 -35.15 ;
    END
  END dout[56]
  PIN dout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.12 -35.47 216.44 -35.15 ;
    END
  END dout[57]
  PIN dout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.24 -35.475 227.56 -35.145 ;
        RECT 227.26 -35.495 227.54 -35.125 ;
    END
  END dout[58]
  PIN dout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.5 -35.47 228.82 -35.15 ;
    END
  END dout[59]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.42 -35.47 22.74 -35.15 ;
    END
  END dout[5]
  PIN dout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.76 -35.47 230.08 -35.15 ;
    END
  END dout[60]
  PIN dout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.02 -35.47 231.34 -35.15 ;
    END
  END dout[61]
  PIN dout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.14 -35.475 242.46 -35.145 ;
        RECT 242.16 -35.495 242.44 -35.125 ;
    END
  END dout[62]
  PIN dout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.4 -35.47 243.72 -35.15 ;
    END
  END dout[63]
  PIN dout[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.66 -35.47 244.98 -35.15 ;
    END
  END dout[64]
  PIN dout[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.92 -35.47 246.24 -35.15 ;
    END
  END dout[65]
  PIN dout[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.04 -35.475 257.36 -35.145 ;
        RECT 257.06 -35.495 257.34 -35.125 ;
    END
  END dout[66]
  PIN dout[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.3 -35.47 258.62 -35.15 ;
    END
  END dout[67]
  PIN dout[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.56 -35.47 259.88 -35.15 ;
    END
  END dout[68]
  PIN dout[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.82 -35.47 261.14 -35.15 ;
    END
  END dout[69]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.54 -35.475 33.86 -35.145 ;
        RECT 33.56 -35.495 33.84 -35.125 ;
    END
  END dout[6]
  PIN dout[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.94 -35.475 272.26 -35.145 ;
        RECT 271.96 -35.495 272.24 -35.125 ;
    END
  END dout[70]
  PIN dout[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.2 -35.47 273.52 -35.15 ;
    END
  END dout[71]
  PIN dout[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.46 -35.47 274.78 -35.15 ;
    END
  END dout[72]
  PIN dout[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.72 -35.47 276.04 -35.15 ;
    END
  END dout[73]
  PIN dout[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.84 -35.475 287.16 -35.145 ;
        RECT 286.86 -35.495 287.14 -35.125 ;
    END
  END dout[74]
  PIN dout[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.1 -35.47 288.42 -35.15 ;
    END
  END dout[75]
  PIN dout[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.36 -35.47 289.68 -35.15 ;
    END
  END dout[76]
  PIN dout[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.62 -35.47 290.94 -35.15 ;
    END
  END dout[77]
  PIN dout[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.74 -35.475 302.06 -35.145 ;
        RECT 301.76 -35.495 302.04 -35.125 ;
    END
  END dout[78]
  PIN dout[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303 -35.47 303.32 -35.15 ;
    END
  END dout[79]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.8 -35.47 35.12 -35.15 ;
    END
  END dout[7]
  PIN dout[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.26 -35.47 304.58 -35.15 ;
    END
  END dout[80]
  PIN dout[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.52 -35.47 305.84 -35.15 ;
    END
  END dout[81]
  PIN dout[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.64 -35.475 316.96 -35.145 ;
        RECT 316.66 -35.495 316.94 -35.125 ;
    END
  END dout[82]
  PIN dout[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.9 -35.47 318.22 -35.15 ;
    END
  END dout[83]
  PIN dout[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.16 -35.47 319.48 -35.15 ;
    END
  END dout[84]
  PIN dout[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.42 -35.47 320.74 -35.15 ;
    END
  END dout[85]
  PIN dout[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.54 -35.475 331.86 -35.145 ;
        RECT 331.56 -35.495 331.84 -35.125 ;
    END
  END dout[86]
  PIN dout[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.8 -35.47 333.12 -35.15 ;
    END
  END dout[87]
  PIN dout[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.06 -35.47 334.38 -35.15 ;
    END
  END dout[88]
  PIN dout[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.32 -35.47 335.64 -35.15 ;
    END
  END dout[89]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.06 -35.47 36.38 -35.15 ;
    END
  END dout[8]
  PIN dout[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.44 -35.475 346.76 -35.145 ;
        RECT 346.46 -35.495 346.74 -35.125 ;
    END
  END dout[90]
  PIN dout[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.7 -35.47 348.02 -35.15 ;
    END
  END dout[91]
  PIN dout[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.96 -35.47 349.28 -35.15 ;
    END
  END dout[92]
  PIN dout[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.22 -35.47 350.54 -35.15 ;
    END
  END dout[93]
  PIN dout[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.34 -35.475 361.66 -35.145 ;
        RECT 361.36 -35.495 361.64 -35.125 ;
    END
  END dout[94]
  PIN dout[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.6 -35.47 362.92 -35.15 ;
    END
  END dout[95]
  PIN dout[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.86 -35.47 364.18 -35.15 ;
    END
  END dout[96]
  PIN dout[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.12 -35.47 365.44 -35.15 ;
    END
  END dout[97]
  PIN dout[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.24 -35.475 376.56 -35.145 ;
        RECT 376.26 -35.495 376.54 -35.125 ;
    END
  END dout[98]
  PIN dout[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.5 -35.47 377.82 -35.15 ;
    END
  END dout[99]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.32 -35.47 37.64 -35.15 ;
    END
  END dout[9]
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -1.36 -22.025 -1.03 -21.695 ;
    END
  END b
  PIN reset_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -1.36 -24.725 -1.03 -24.395 ;
    END
  END reset_b
  OBS
    LAYER met1 ;
      RECT 946.22 -35.47 949.06 -35.15 ;
      RECT 930.06 -35.47 934.79 -35.15 ;
      RECT 915.16 -35.47 919.89 -35.15 ;
      RECT 900.26 -35.47 904.99 -35.15 ;
      RECT 885.36 -35.47 890.09 -35.15 ;
      RECT 870.46 -35.47 875.19 -35.15 ;
      RECT 855.56 -35.47 860.29 -35.15 ;
      RECT 840.66 -35.47 845.39 -35.15 ;
      RECT 825.76 -35.47 830.49 -35.15 ;
      RECT 810.86 -35.47 815.59 -35.15 ;
      RECT 795.96 -35.47 800.69 -35.15 ;
      RECT 781.06 -35.47 785.79 -35.15 ;
      RECT 766.16 -35.47 770.89 -35.15 ;
      RECT 751.26 -35.47 755.99 -35.15 ;
      RECT 736.36 -35.47 741.09 -35.15 ;
      RECT 721.46 -35.47 726.19 -35.15 ;
      RECT 706.56 -35.47 711.29 -35.15 ;
      RECT 691.66 -35.47 696.39 -35.15 ;
      RECT 676.76 -35.47 681.49 -35.15 ;
      RECT 661.86 -35.47 666.59 -35.15 ;
      RECT 646.96 -35.47 651.69 -35.15 ;
      RECT 632.06 -35.47 636.79 -35.15 ;
      RECT 617.16 -35.47 621.89 -35.15 ;
      RECT 602.26 -35.47 606.99 -35.15 ;
      RECT 587.36 -35.47 592.09 -35.15 ;
      RECT 572.46 -35.47 577.19 -35.15 ;
      RECT 557.56 -35.47 562.29 -35.15 ;
      RECT 542.66 -35.47 547.39 -35.15 ;
      RECT 527.76 -35.47 532.49 -35.15 ;
      RECT 512.86 -35.47 517.59 -35.15 ;
      RECT 497.96 -35.47 502.69 -35.15 ;
      RECT 483.06 -35.47 487.79 -35.15 ;
      RECT 468.16 -35.47 472.89 -35.15 ;
      RECT 453.26 -35.47 457.99 -35.15 ;
      RECT 438.36 -35.47 443.09 -35.15 ;
      RECT 423.46 -35.47 428.19 -35.15 ;
      RECT 408.56 -35.47 413.29 -35.15 ;
      RECT 393.66 -35.47 398.39 -35.15 ;
      RECT 378.76 -35.47 383.49 -35.15 ;
      RECT 363.86 -35.47 368.59 -35.15 ;
      RECT 348.96 -35.47 353.69 -35.15 ;
      RECT 334.06 -35.47 338.79 -35.15 ;
      RECT 319.16 -35.47 323.89 -35.15 ;
      RECT 304.26 -35.47 308.99 -35.15 ;
      RECT 289.36 -35.47 294.09 -35.15 ;
      RECT 274.46 -35.47 279.19 -35.15 ;
      RECT 259.56 -35.47 264.29 -35.15 ;
      RECT 244.66 -35.47 249.39 -35.15 ;
      RECT 229.76 -35.47 234.49 -35.15 ;
      RECT 214.86 -35.47 219.59 -35.15 ;
      RECT 199.96 -35.47 204.69 -35.15 ;
      RECT 185.06 -35.47 189.79 -35.15 ;
      RECT 170.16 -35.47 174.89 -35.15 ;
      RECT 155.26 -35.47 159.99 -35.15 ;
      RECT 140.36 -35.47 145.09 -35.15 ;
      RECT 125.46 -35.47 130.19 -35.15 ;
      RECT 110.56 -35.47 115.29 -35.15 ;
      RECT 95.66 -35.47 100.39 -35.15 ;
      RECT 80.76 -35.47 85.49 -35.15 ;
      RECT 65.86 -35.47 70.59 -35.15 ;
      RECT 50.96 -35.47 55.69 -35.15 ;
      RECT 36.06 -35.47 40.79 -35.15 ;
      RECT 21.16 -35.47 25.89 -35.15 ;
      RECT 7.52 -35.47 10.36 -35.15 ;
    LAYER met1 SPACING 0.14 ;
      RECT -1.525 -35.545 954.885 2.225 ;
    LAYER met2 ;
      RECT 954.56 -35.52 954.88 2.2 ;
      RECT 954.58 -35.545 954.86 2.2 ;
      RECT 953.9 -35.52 954.18 2.225 ;
      RECT 953.88 -35.52 954.2 2.2 ;
      RECT 953.2 -35.52 953.52 2.2 ;
      RECT 953.22 -35.545 953.5 2.2 ;
      RECT 952.54 -35.52 952.82 2.225 ;
      RECT 952.52 -35.52 952.84 2.2 ;
      RECT 951.84 -35.52 952.16 2.2 ;
      RECT 951.86 -35.545 952.14 2.2 ;
      RECT 951.18 -35.52 951.46 2.225 ;
      RECT 951.16 -35.52 951.48 2.2 ;
      RECT 950.48 -35.52 950.8 2.2 ;
      RECT 950.5 -35.545 950.78 2.2 ;
      RECT 949.82 -35.52 950.1 2.225 ;
      RECT 949.8 -35.52 950.12 2.2 ;
      RECT 948.46 -20.56 948.74 2.225 ;
      RECT 948.44 -20.56 948.76 2.2 ;
      RECT 948.11 -35.475 948.43 -25.07 ;
      RECT 948.13 -35.495 948.41 -25.07 ;
      RECT 947.1 -35.52 947.38 2.225 ;
      RECT 947.08 -35.52 947.4 2.2 ;
      RECT 945.74 -34.16 946.02 2.225 ;
      RECT 945.72 -34.16 946.04 2.2 ;
      RECT 944.38 -18.52 944.66 2.225 ;
      RECT 944.36 -18.52 944.68 2.2 ;
      RECT 943.68 -35.52 944 -23.64 ;
      RECT 943.7 -35.545 943.98 -23.64 ;
      RECT 943.02 -21.92 943.3 2.225 ;
      RECT 943 -21.92 943.32 2.2 ;
      RECT 942.32 -35.52 942.64 -25 ;
      RECT 942.34 -35.545 942.62 -25 ;
      RECT 941.66 -18.52 941.94 2.225 ;
      RECT 941.64 -18.52 941.96 2.2 ;
      RECT 940.96 -35.52 941.28 -25.68 ;
      RECT 940.98 -35.545 941.26 -25.68 ;
      RECT 940.3 -35.52 940.58 2.225 ;
      RECT 940.28 -35.52 940.6 2.2 ;
      RECT 939.6 -35.52 939.92 2.2 ;
      RECT 939.62 -35.545 939.9 2.2 ;
      RECT 938.94 -35.52 939.22 2.225 ;
      RECT 938.92 -35.52 939.24 2.2 ;
      RECT 938.24 -35.52 938.56 2.2 ;
      RECT 938.26 -35.545 938.54 2.2 ;
      RECT 937.58 -35.52 937.86 2.225 ;
      RECT 937.56 -35.52 937.88 2.2 ;
      RECT 936.88 -35.52 937.2 2.2 ;
      RECT 936.9 -35.545 937.18 2.2 ;
      RECT 936.22 -35.52 936.5 2.225 ;
      RECT 936.2 -35.52 936.52 2.2 ;
      RECT 935.52 -35.52 935.84 2.2 ;
      RECT 935.54 -35.545 935.82 2.2 ;
      RECT 934.86 -24.64 935.14 2.225 ;
      RECT 934.84 -24.64 935.16 2.2 ;
      RECT 933.84 -35.475 934.16 -30.11 ;
      RECT 933.86 -35.495 934.14 -30.11 ;
      RECT 933.5 -20.56 933.78 2.225 ;
      RECT 933.48 -20.56 933.8 2.2 ;
      RECT 932.14 -35.52 932.42 2.225 ;
      RECT 932.12 -35.52 932.44 2.2 ;
      RECT 930.78 -25.32 931.06 2.225 ;
      RECT 930.76 -25.32 931.08 2.2 ;
      RECT 929.42 -17.16 929.7 2.225 ;
      RECT 929.4 -17.16 929.72 2.2 ;
      RECT 928.06 -21.92 928.34 2.225 ;
      RECT 928.04 -21.92 928.36 2.2 ;
      RECT 926.7 -18.52 926.98 2.225 ;
      RECT 926.68 -18.52 927 2.2 ;
      RECT 926 -35.52 926.32 -31.12 ;
      RECT 926.02 -35.545 926.3 -31.12 ;
      RECT 925.34 -35.52 925.62 2.225 ;
      RECT 925.32 -35.52 925.64 2.2 ;
      RECT 924.64 -35.52 924.96 2.2 ;
      RECT 924.66 -35.545 924.94 2.2 ;
      RECT 923.98 -35.52 924.26 2.225 ;
      RECT 923.96 -35.52 924.28 2.2 ;
      RECT 923.28 -35.52 923.6 2.2 ;
      RECT 923.3 -35.545 923.58 2.2 ;
      RECT 922.62 -35.52 922.9 2.225 ;
      RECT 922.6 -35.52 922.92 2.2 ;
      RECT 921.92 -35.52 922.24 2.2 ;
      RECT 921.94 -35.545 922.22 2.2 ;
      RECT 921.26 -35.52 921.54 2.225 ;
      RECT 921.24 -35.52 921.56 2.2 ;
      RECT 920.56 -35.52 920.88 2.2 ;
      RECT 920.58 -35.545 920.86 2.2 ;
      RECT 919.9 -24.64 920.18 2.225 ;
      RECT 919.88 -24.64 920.2 2.2 ;
      RECT 918.94 -35.475 919.26 -30.11 ;
      RECT 918.96 -35.495 919.24 -30.11 ;
      RECT 918.54 -20.56 918.82 2.225 ;
      RECT 918.52 -20.56 918.84 2.2 ;
      RECT 917.18 -35.52 917.46 2.225 ;
      RECT 917.16 -35.52 917.48 2.2 ;
      RECT 915.82 -17.16 916.1 2.225 ;
      RECT 915.8 -17.16 916.12 2.2 ;
      RECT 914.46 -17.84 914.74 2.225 ;
      RECT 914.44 -17.84 914.76 2.2 ;
      RECT 913.1 -21.92 913.38 2.225 ;
      RECT 913.08 -21.92 913.4 2.2 ;
      RECT 911.74 -18.52 912.02 2.225 ;
      RECT 911.72 -18.52 912.04 2.2 ;
      RECT 911.04 -35.52 911.36 -31.12 ;
      RECT 911.06 -35.545 911.34 -31.12 ;
      RECT 910.38 -35.52 910.66 2.225 ;
      RECT 910.36 -35.52 910.68 2.2 ;
      RECT 909.68 -35.52 910 2.2 ;
      RECT 909.7 -35.545 909.98 2.2 ;
      RECT 909.02 -35.52 909.3 2.225 ;
      RECT 909 -35.52 909.32 2.2 ;
      RECT 908.32 -35.52 908.64 2.2 ;
      RECT 908.34 -35.545 908.62 2.2 ;
      RECT 907.66 -35.52 907.94 2.225 ;
      RECT 907.64 -35.52 907.96 2.2 ;
      RECT 906.96 -35.52 907.28 2.2 ;
      RECT 906.98 -35.545 907.26 2.2 ;
      RECT 906.3 -35.52 906.58 2.225 ;
      RECT 906.28 -35.52 906.6 2.2 ;
      RECT 905.6 -35.52 905.92 2.2 ;
      RECT 905.62 -35.545 905.9 2.2 ;
      RECT 904.94 -24.64 905.22 2.225 ;
      RECT 904.92 -24.64 905.24 2.2 ;
      RECT 904.04 -35.475 904.36 -30.11 ;
      RECT 904.06 -35.495 904.34 -30.11 ;
      RECT 903.58 -20.56 903.86 2.225 ;
      RECT 903.56 -20.56 903.88 2.2 ;
      RECT 902.22 -35.52 902.5 2.225 ;
      RECT 902.2 -35.52 902.52 2.2 ;
      RECT 900.86 -17.16 901.14 2.225 ;
      RECT 900.84 -17.16 901.16 2.2 ;
      RECT 899.5 -17.84 899.78 2.225 ;
      RECT 899.48 -17.84 899.8 2.2 ;
      RECT 898.14 -21.92 898.42 2.225 ;
      RECT 898.12 -21.92 898.44 2.2 ;
      RECT 896.78 -18.52 897.06 2.225 ;
      RECT 896.76 -18.52 897.08 2.2 ;
      RECT 896.08 -35.52 896.4 -31.12 ;
      RECT 896.1 -35.545 896.38 -31.12 ;
      RECT 895.42 -35.52 895.7 2.225 ;
      RECT 895.4 -35.52 895.72 2.2 ;
      RECT 894.72 -35.52 895.04 2.2 ;
      RECT 894.74 -35.545 895.02 2.2 ;
      RECT 894.06 -35.52 894.34 2.225 ;
      RECT 894.04 -35.52 894.36 2.2 ;
      RECT 893.36 -35.52 893.68 2.2 ;
      RECT 893.38 -35.545 893.66 2.2 ;
      RECT 892.7 -35.52 892.98 2.225 ;
      RECT 892.68 -35.52 893 2.2 ;
      RECT 892 -35.52 892.32 2.2 ;
      RECT 892.02 -35.545 892.3 2.2 ;
      RECT 891.34 -35.52 891.62 2.225 ;
      RECT 891.32 -35.52 891.64 2.2 ;
      RECT 890.64 -35.52 890.96 2.2 ;
      RECT 890.66 -35.545 890.94 2.2 ;
      RECT 889.98 -24.64 890.26 2.225 ;
      RECT 889.96 -24.64 890.28 2.2 ;
      RECT 889.14 -35.475 889.46 -30.11 ;
      RECT 889.16 -35.495 889.44 -30.11 ;
      RECT 888.62 -20.56 888.9 2.225 ;
      RECT 888.6 -20.56 888.92 2.2 ;
      RECT 887.26 -25.32 887.54 2.225 ;
      RECT 887.24 -25.32 887.56 2.2 ;
      RECT 885.9 -17.16 886.18 2.225 ;
      RECT 885.88 -17.16 886.2 2.2 ;
      RECT 884.54 -17.84 884.82 2.225 ;
      RECT 884.52 -17.84 884.84 2.2 ;
      RECT 883.18 -21.92 883.46 2.225 ;
      RECT 883.16 -21.92 883.48 2.2 ;
      RECT 881.82 -18.52 882.1 2.225 ;
      RECT 881.8 -18.52 882.12 2.2 ;
      RECT 881.12 -35.52 881.44 -31.12 ;
      RECT 881.14 -35.545 881.42 -31.12 ;
      RECT 880.46 -35.52 880.74 2.225 ;
      RECT 880.44 -35.52 880.76 2.2 ;
      RECT 879.76 -35.52 880.08 2.2 ;
      RECT 879.78 -35.545 880.06 2.2 ;
      RECT 879.1 -35.52 879.38 2.225 ;
      RECT 879.08 -35.52 879.4 2.2 ;
      RECT 878.4 -35.52 878.72 2.2 ;
      RECT 878.42 -35.545 878.7 2.2 ;
      RECT 877.74 -35.52 878.02 2.225 ;
      RECT 877.72 -35.52 878.04 2.2 ;
      RECT 877.04 -35.52 877.36 2.2 ;
      RECT 877.06 -35.545 877.34 2.2 ;
      RECT 876.38 -35.52 876.66 2.225 ;
      RECT 876.36 -35.52 876.68 2.2 ;
      RECT 875.68 -35.52 876 2.2 ;
      RECT 875.7 -35.545 875.98 2.2 ;
      RECT 875.02 -24.64 875.3 2.225 ;
      RECT 875 -24.64 875.32 2.2 ;
      RECT 874.24 -35.475 874.56 -30.11 ;
      RECT 874.26 -35.495 874.54 -30.11 ;
      RECT 873.66 -20.56 873.94 2.225 ;
      RECT 873.64 -20.56 873.96 2.2 ;
      RECT 872.3 -25.32 872.58 2.225 ;
      RECT 872.28 -25.32 872.6 2.2 ;
      RECT 870.94 -17.16 871.22 2.225 ;
      RECT 870.92 -17.16 871.24 2.2 ;
      RECT 869.58 -17.84 869.86 2.225 ;
      RECT 869.56 -17.84 869.88 2.2 ;
      RECT 868.22 -21.92 868.5 2.225 ;
      RECT 868.2 -21.92 868.52 2.2 ;
      RECT 866.86 -18.52 867.14 2.225 ;
      RECT 866.84 -18.52 867.16 2.2 ;
      RECT 866.16 -35.52 866.48 -31.12 ;
      RECT 866.18 -35.545 866.46 -31.12 ;
      RECT 865.5 -35.52 865.78 2.225 ;
      RECT 865.48 -35.52 865.8 2.2 ;
      RECT 864.8 -35.52 865.12 2.2 ;
      RECT 864.82 -35.545 865.1 2.2 ;
      RECT 864.14 -35.52 864.42 2.225 ;
      RECT 864.12 -35.52 864.44 2.2 ;
      RECT 863.44 -35.52 863.76 2.2 ;
      RECT 863.46 -35.545 863.74 2.2 ;
      RECT 862.78 -35.52 863.06 2.225 ;
      RECT 862.76 -35.52 863.08 2.2 ;
      RECT 862.08 -35.52 862.4 2.2 ;
      RECT 862.1 -35.545 862.38 2.2 ;
      RECT 861.42 -35.52 861.7 2.225 ;
      RECT 861.4 -35.52 861.72 2.2 ;
      RECT 860.72 -35.52 861.04 2.2 ;
      RECT 860.74 -35.545 861.02 2.2 ;
      RECT 860.06 -24.64 860.34 2.225 ;
      RECT 860.04 -24.64 860.36 2.2 ;
      RECT 859.34 -35.475 859.66 -30.11 ;
      RECT 859.36 -35.495 859.64 -30.11 ;
      RECT 858.7 -20.56 858.98 2.225 ;
      RECT 858.68 -20.56 859 2.2 ;
      RECT 857.34 -25.32 857.62 2.225 ;
      RECT 857.32 -25.32 857.64 2.2 ;
      RECT 855.98 -17.16 856.26 2.225 ;
      RECT 855.96 -17.16 856.28 2.2 ;
      RECT 854.62 -17.84 854.9 2.225 ;
      RECT 854.6 -17.84 854.92 2.2 ;
      RECT 853.26 -21.92 853.54 2.225 ;
      RECT 853.24 -21.92 853.56 2.2 ;
      RECT 851.9 -18.52 852.18 2.225 ;
      RECT 851.88 -18.52 852.2 2.2 ;
      RECT 851.2 -35.52 851.52 -31.12 ;
      RECT 851.22 -35.545 851.5 -31.12 ;
      RECT 850.54 -35.52 850.82 2.225 ;
      RECT 850.52 -35.52 850.84 2.2 ;
      RECT 849.84 -35.52 850.16 2.2 ;
      RECT 849.86 -35.545 850.14 2.2 ;
      RECT 849.18 -35.52 849.46 2.225 ;
      RECT 849.16 -35.52 849.48 2.2 ;
      RECT 848.48 -35.52 848.8 2.2 ;
      RECT 848.5 -35.545 848.78 2.2 ;
      RECT 847.82 -35.52 848.1 2.225 ;
      RECT 847.8 -35.52 848.12 2.2 ;
      RECT 847.12 -35.52 847.44 2.2 ;
      RECT 847.14 -35.545 847.42 2.2 ;
      RECT 846.46 -35.52 846.74 2.225 ;
      RECT 846.44 -35.52 846.76 2.2 ;
      RECT 845.76 -35.52 846.08 2.2 ;
      RECT 845.78 -35.545 846.06 2.2 ;
      RECT 845.1 -20.56 845.38 2.225 ;
      RECT 845.08 -20.56 845.4 2.2 ;
      RECT 844.44 -35.475 844.76 -30.11 ;
      RECT 844.46 -35.495 844.74 -30.11 ;
      RECT 843.74 -21.24 844.02 2.225 ;
      RECT 843.72 -21.24 844.04 2.2 ;
      RECT 842.38 -25.32 842.66 2.225 ;
      RECT 842.36 -25.32 842.68 2.2 ;
      RECT 841.02 -17.16 841.3 2.225 ;
      RECT 841 -17.16 841.32 2.2 ;
      RECT 839.66 -17.84 839.94 2.225 ;
      RECT 839.64 -17.84 839.96 2.2 ;
      RECT 838.3 -21.92 838.58 2.225 ;
      RECT 838.28 -21.92 838.6 2.2 ;
      RECT 836.94 -18.52 837.22 2.225 ;
      RECT 836.92 -18.52 837.24 2.2 ;
      RECT 836.24 -35.52 836.56 -31.12 ;
      RECT 836.26 -35.545 836.54 -31.12 ;
      RECT 835.58 -35.52 835.86 2.225 ;
      RECT 835.56 -35.52 835.88 2.2 ;
      RECT 834.88 -35.52 835.2 2.2 ;
      RECT 834.9 -35.545 835.18 2.2 ;
      RECT 834.22 -35.52 834.5 2.225 ;
      RECT 834.2 -35.52 834.52 2.2 ;
      RECT 833.52 -35.52 833.84 2.2 ;
      RECT 833.54 -35.545 833.82 2.2 ;
      RECT 832.86 -35.52 833.14 2.225 ;
      RECT 832.84 -35.52 833.16 2.2 ;
      RECT 832.16 -35.52 832.48 2.2 ;
      RECT 832.18 -35.545 832.46 2.2 ;
      RECT 831.5 -35.52 831.78 2.225 ;
      RECT 831.48 -35.52 831.8 2.2 ;
      RECT 830.14 -20.56 830.42 2.225 ;
      RECT 830.12 -20.56 830.44 2.2 ;
      RECT 829.54 -35.475 829.86 -30.11 ;
      RECT 829.56 -35.495 829.84 -30.11 ;
      RECT 828.78 -21.24 829.06 2.225 ;
      RECT 828.76 -21.24 829.08 2.2 ;
      RECT 827.42 -25.32 827.7 2.225 ;
      RECT 827.4 -25.32 827.72 2.2 ;
      RECT 826.06 -17.16 826.34 2.225 ;
      RECT 826.04 -17.16 826.36 2.2 ;
      RECT 824.7 -17.84 824.98 2.225 ;
      RECT 824.68 -17.84 825 2.2 ;
      RECT 823.34 -21.92 823.62 2.225 ;
      RECT 823.32 -21.92 823.64 2.2 ;
      RECT 821.98 -18.52 822.26 2.225 ;
      RECT 821.96 -18.52 822.28 2.2 ;
      RECT 821.28 -35.52 821.6 -31.12 ;
      RECT 821.3 -35.545 821.58 -31.12 ;
      RECT 820.62 -35.52 820.9 2.225 ;
      RECT 820.6 -35.52 820.92 2.2 ;
      RECT 819.92 -35.52 820.24 2.2 ;
      RECT 819.94 -35.545 820.22 2.2 ;
      RECT 819.26 -35.52 819.54 2.225 ;
      RECT 819.24 -35.52 819.56 2.2 ;
      RECT 818.56 -35.52 818.88 2.2 ;
      RECT 818.58 -35.545 818.86 2.2 ;
      RECT 817.9 -35.52 818.18 2.225 ;
      RECT 817.88 -35.52 818.2 2.2 ;
      RECT 817.2 -35.52 817.52 2.2 ;
      RECT 817.22 -35.545 817.5 2.2 ;
      RECT 816.54 -35.52 816.82 2.225 ;
      RECT 816.52 -35.52 816.84 2.2 ;
      RECT 815.18 -20.56 815.46 2.225 ;
      RECT 815.16 -20.56 815.48 2.2 ;
      RECT 814.64 -35.475 814.96 -30.11 ;
      RECT 814.66 -35.495 814.94 -30.11 ;
      RECT 813.82 -21.24 814.1 2.225 ;
      RECT 813.8 -21.24 814.12 2.2 ;
      RECT 812.46 -25.32 812.74 2.225 ;
      RECT 812.44 -25.32 812.76 2.2 ;
      RECT 811.1 -17.16 811.38 2.225 ;
      RECT 811.08 -17.16 811.4 2.2 ;
      RECT 809.74 -17.84 810.02 2.225 ;
      RECT 809.72 -17.84 810.04 2.2 ;
      RECT 808.38 -18.52 808.66 2.225 ;
      RECT 808.36 -18.52 808.68 2.2 ;
      RECT 807.02 -21.24 807.3 2.225 ;
      RECT 807 -21.24 807.32 2.2 ;
      RECT 806.32 -35.52 806.64 -31.12 ;
      RECT 806.34 -35.545 806.62 -31.12 ;
      RECT 805.66 -35.52 805.94 2.225 ;
      RECT 805.64 -35.52 805.96 2.2 ;
      RECT 804.96 -35.52 805.28 2.2 ;
      RECT 804.98 -35.545 805.26 2.2 ;
      RECT 804.3 -35.52 804.58 2.225 ;
      RECT 804.28 -35.52 804.6 2.2 ;
      RECT 803.6 -35.52 803.92 2.2 ;
      RECT 803.62 -35.545 803.9 2.2 ;
      RECT 802.94 -35.52 803.22 2.225 ;
      RECT 802.92 -35.52 803.24 2.2 ;
      RECT 802.24 -35.52 802.56 2.2 ;
      RECT 802.26 -35.545 802.54 2.2 ;
      RECT 801.58 -35.52 801.86 2.225 ;
      RECT 801.56 -35.52 801.88 2.2 ;
      RECT 800.22 -20.56 800.5 2.225 ;
      RECT 800.2 -20.56 800.52 2.2 ;
      RECT 799.74 -35.475 800.06 -30.11 ;
      RECT 799.76 -35.495 800.04 -30.11 ;
      RECT 798.86 -21.24 799.14 2.225 ;
      RECT 798.84 -21.24 799.16 2.2 ;
      RECT 797.5 -25.32 797.78 2.225 ;
      RECT 797.48 -25.32 797.8 2.2 ;
      RECT 796.14 -17.16 796.42 2.225 ;
      RECT 796.12 -17.16 796.44 2.2 ;
      RECT 794.78 -17.84 795.06 2.225 ;
      RECT 794.76 -17.84 795.08 2.2 ;
      RECT 793.42 -18.52 793.7 2.225 ;
      RECT 793.4 -18.52 793.72 2.2 ;
      RECT 792.72 -35.52 793.04 -31.12 ;
      RECT 792.74 -35.545 793.02 -31.12 ;
      RECT 792.06 -21.24 792.34 2.225 ;
      RECT 792.04 -21.24 792.36 2.2 ;
      RECT 791.36 -35.52 791.68 2.2 ;
      RECT 791.38 -35.545 791.66 2.2 ;
      RECT 790.7 -35.52 790.98 2.225 ;
      RECT 790.68 -35.52 791 2.2 ;
      RECT 790 -35.52 790.32 2.2 ;
      RECT 790.02 -35.545 790.3 2.2 ;
      RECT 789.34 -35.52 789.62 2.225 ;
      RECT 789.32 -35.52 789.64 2.2 ;
      RECT 788.64 -35.52 788.96 2.2 ;
      RECT 788.66 -35.545 788.94 2.2 ;
      RECT 787.98 -35.52 788.26 2.225 ;
      RECT 787.96 -35.52 788.28 2.2 ;
      RECT 787.28 -35.52 787.6 2.2 ;
      RECT 787.3 -35.545 787.58 2.2 ;
      RECT 786.62 -35.52 786.9 2.225 ;
      RECT 786.6 -35.52 786.92 2.2 ;
      RECT 785.26 -20.56 785.54 2.225 ;
      RECT 785.24 -20.56 785.56 2.2 ;
      RECT 784.84 -35.475 785.16 -30.11 ;
      RECT 784.86 -35.495 785.14 -30.11 ;
      RECT 783.9 -21.24 784.18 2.225 ;
      RECT 783.88 -21.24 784.2 2.2 ;
      RECT 782.54 -25.32 782.82 2.225 ;
      RECT 782.52 -25.32 782.84 2.2 ;
      RECT 781.18 -17.16 781.46 2.225 ;
      RECT 781.16 -17.16 781.48 2.2 ;
      RECT 779.82 -17.84 780.1 2.225 ;
      RECT 779.8 -17.84 780.12 2.2 ;
      RECT 778.46 -18.52 778.74 2.225 ;
      RECT 778.44 -18.52 778.76 2.2 ;
      RECT 777.76 -35.52 778.08 -31.12 ;
      RECT 777.78 -35.545 778.06 -31.12 ;
      RECT 777.1 -21.24 777.38 2.225 ;
      RECT 777.08 -21.24 777.4 2.2 ;
      RECT 776.4 -35.52 776.72 2.2 ;
      RECT 776.42 -35.545 776.7 2.2 ;
      RECT 775.74 -35.52 776.02 2.225 ;
      RECT 775.72 -35.52 776.04 2.2 ;
      RECT 775.04 -35.52 775.36 2.2 ;
      RECT 775.06 -35.545 775.34 2.2 ;
      RECT 774.38 -35.52 774.66 2.225 ;
      RECT 774.36 -35.52 774.68 2.2 ;
      RECT 773.68 -35.52 774 2.2 ;
      RECT 773.7 -35.545 773.98 2.2 ;
      RECT 773.02 -35.52 773.3 2.225 ;
      RECT 773 -35.52 773.32 2.2 ;
      RECT 772.32 -35.52 772.64 2.2 ;
      RECT 772.34 -35.545 772.62 2.2 ;
      RECT 771.66 -35.52 771.94 2.225 ;
      RECT 771.64 -35.52 771.96 2.2 ;
      RECT 770.3 -20.56 770.58 2.225 ;
      RECT 770.28 -20.56 770.6 2.2 ;
      RECT 769.94 -35.475 770.26 -30.11 ;
      RECT 769.96 -35.495 770.24 -30.11 ;
      RECT 768.94 -21.24 769.22 2.225 ;
      RECT 768.92 -21.24 769.24 2.2 ;
      RECT 767.58 -25.32 767.86 2.225 ;
      RECT 767.56 -25.32 767.88 2.2 ;
      RECT 766.22 -17.16 766.5 2.225 ;
      RECT 766.2 -17.16 766.52 2.2 ;
      RECT 764.86 -18.52 765.14 2.225 ;
      RECT 764.84 -18.52 765.16 2.2 ;
      RECT 763.5 -18.52 763.78 2.225 ;
      RECT 763.48 -18.52 763.8 2.2 ;
      RECT 762.8 -35.52 763.12 -31.12 ;
      RECT 762.82 -35.545 763.1 -31.12 ;
      RECT 762.14 -21.24 762.42 2.225 ;
      RECT 762.12 -21.24 762.44 2.2 ;
      RECT 761.44 -35.52 761.76 2.2 ;
      RECT 761.46 -35.545 761.74 2.2 ;
      RECT 760.78 -35.52 761.06 2.225 ;
      RECT 760.76 -35.52 761.08 2.2 ;
      RECT 760.08 -35.52 760.4 2.2 ;
      RECT 760.1 -35.545 760.38 2.2 ;
      RECT 759.42 -35.52 759.7 2.225 ;
      RECT 759.4 -35.52 759.72 2.2 ;
      RECT 758.72 -35.52 759.04 2.2 ;
      RECT 758.74 -35.545 759.02 2.2 ;
      RECT 758.06 -35.52 758.34 2.225 ;
      RECT 758.04 -35.52 758.36 2.2 ;
      RECT 757.36 -35.52 757.68 2.2 ;
      RECT 757.38 -35.545 757.66 2.2 ;
      RECT 756.7 -35.52 756.98 2.225 ;
      RECT 756.68 -35.52 757 2.2 ;
      RECT 755.34 -20.56 755.62 2.225 ;
      RECT 755.32 -20.56 755.64 2.2 ;
      RECT 755.04 -35.475 755.36 -30.11 ;
      RECT 755.06 -35.495 755.34 -30.11 ;
      RECT 753.98 -21.24 754.26 2.225 ;
      RECT 753.96 -21.24 754.28 2.2 ;
      RECT 752.62 -25.32 752.9 2.225 ;
      RECT 752.6 -25.32 752.92 2.2 ;
      RECT 751.26 -17.16 751.54 2.225 ;
      RECT 751.24 -17.16 751.56 2.2 ;
      RECT 749.9 -18.52 750.18 2.225 ;
      RECT 749.88 -18.52 750.2 2.2 ;
      RECT 748.54 -18.52 748.82 2.225 ;
      RECT 748.52 -18.52 748.84 2.2 ;
      RECT 747.84 -35.52 748.16 -31.12 ;
      RECT 747.86 -35.545 748.14 -31.12 ;
      RECT 747.18 -21.24 747.46 2.225 ;
      RECT 747.16 -21.24 747.48 2.2 ;
      RECT 746.48 -35.52 746.8 2.2 ;
      RECT 746.5 -35.545 746.78 2.2 ;
      RECT 745.82 -35.52 746.1 2.225 ;
      RECT 745.8 -35.52 746.12 2.2 ;
      RECT 745.12 -35.52 745.44 2.2 ;
      RECT 745.14 -35.545 745.42 2.2 ;
      RECT 744.46 -35.52 744.74 2.225 ;
      RECT 744.44 -35.52 744.76 2.2 ;
      RECT 743.76 -35.52 744.08 2.2 ;
      RECT 743.78 -35.545 744.06 2.2 ;
      RECT 743.1 -35.52 743.38 2.225 ;
      RECT 743.08 -35.52 743.4 2.2 ;
      RECT 742.4 -35.52 742.72 2.2 ;
      RECT 742.42 -35.545 742.7 2.2 ;
      RECT 741.74 -35.52 742.02 2.225 ;
      RECT 741.72 -35.52 742.04 2.2 ;
      RECT 740.38 -20.56 740.66 2.225 ;
      RECT 740.36 -20.56 740.68 2.2 ;
      RECT 740.14 -35.475 740.46 -30.11 ;
      RECT 740.16 -35.495 740.44 -30.11 ;
      RECT 739.02 -21.24 739.3 2.225 ;
      RECT 739 -21.24 739.32 2.2 ;
      RECT 737.66 -25.32 737.94 2.225 ;
      RECT 737.64 -25.32 737.96 2.2 ;
      RECT 736.3 -17.16 736.58 2.225 ;
      RECT 736.28 -17.16 736.6 2.2 ;
      RECT 734.94 -18.52 735.22 2.225 ;
      RECT 734.92 -18.52 735.24 2.2 ;
      RECT 733.58 -18.52 733.86 2.225 ;
      RECT 733.56 -18.52 733.88 2.2 ;
      RECT 732.88 -35.52 733.2 -31.12 ;
      RECT 732.9 -35.545 733.18 -31.12 ;
      RECT 732.22 -21.24 732.5 2.225 ;
      RECT 732.2 -21.24 732.52 2.2 ;
      RECT 731.52 -35.52 731.84 2.2 ;
      RECT 731.54 -35.545 731.82 2.2 ;
      RECT 730.86 -35.52 731.14 2.225 ;
      RECT 730.84 -35.52 731.16 2.2 ;
      RECT 730.16 -35.52 730.48 2.2 ;
      RECT 730.18 -35.545 730.46 2.2 ;
      RECT 729.5 -35.52 729.78 2.225 ;
      RECT 729.48 -35.52 729.8 2.2 ;
      RECT 728.8 -35.52 729.12 2.2 ;
      RECT 728.82 -35.545 729.1 2.2 ;
      RECT 728.14 -35.52 728.42 2.225 ;
      RECT 728.12 -35.52 728.44 2.2 ;
      RECT 727.44 -35.52 727.76 2.2 ;
      RECT 727.46 -35.545 727.74 2.2 ;
      RECT 726.78 -35.52 727.06 2.225 ;
      RECT 726.76 -35.52 727.08 2.2 ;
      RECT 725.42 -20.56 725.7 2.225 ;
      RECT 725.4 -20.56 725.72 2.2 ;
      RECT 725.24 -35.475 725.56 -30.11 ;
      RECT 725.26 -35.495 725.54 -30.11 ;
      RECT 724.06 -21.24 724.34 2.225 ;
      RECT 724.04 -21.24 724.36 2.2 ;
      RECT 722.7 -25.32 722.98 2.225 ;
      RECT 722.68 -25.32 723 2.2 ;
      RECT 721.34 -17.16 721.62 2.225 ;
      RECT 721.32 -17.16 721.64 2.2 ;
      RECT 719.98 -18.52 720.26 2.225 ;
      RECT 719.96 -18.52 720.28 2.2 ;
      RECT 718.62 -18.52 718.9 2.225 ;
      RECT 718.6 -18.52 718.92 2.2 ;
      RECT 717.92 -35.52 718.24 -31.12 ;
      RECT 717.94 -35.545 718.22 -31.12 ;
      RECT 717.26 -21.24 717.54 2.225 ;
      RECT 717.24 -21.24 717.56 2.2 ;
      RECT 716.56 -35.52 716.88 2.2 ;
      RECT 716.58 -35.545 716.86 2.2 ;
      RECT 715.9 -35.52 716.18 2.225 ;
      RECT 715.88 -35.52 716.2 2.2 ;
      RECT 715.2 -35.52 715.52 2.2 ;
      RECT 715.22 -35.545 715.5 2.2 ;
      RECT 714.54 -35.52 714.82 2.225 ;
      RECT 714.52 -35.52 714.84 2.2 ;
      RECT 713.84 -35.52 714.16 2.2 ;
      RECT 713.86 -35.545 714.14 2.2 ;
      RECT 713.18 -35.52 713.46 2.225 ;
      RECT 713.16 -35.52 713.48 2.2 ;
      RECT 712.48 -35.52 712.8 2.2 ;
      RECT 712.5 -35.545 712.78 2.2 ;
      RECT 711.82 -35.52 712.1 2.225 ;
      RECT 711.8 -35.52 712.12 2.2 ;
      RECT 710.46 -20.56 710.74 2.225 ;
      RECT 710.44 -20.56 710.76 2.2 ;
      RECT 710.34 -35.475 710.66 -30.11 ;
      RECT 710.36 -35.495 710.64 -30.11 ;
      RECT 709.1 -21.24 709.38 2.225 ;
      RECT 709.08 -21.24 709.4 2.2 ;
      RECT 707.74 -25.32 708.02 2.225 ;
      RECT 707.72 -25.32 708.04 2.2 ;
      RECT 706.38 -17.16 706.66 2.225 ;
      RECT 706.36 -17.16 706.68 2.2 ;
      RECT 705.02 -18.52 705.3 2.225 ;
      RECT 705 -18.52 705.32 2.2 ;
      RECT 703.66 -18.52 703.94 2.225 ;
      RECT 703.64 -18.52 703.96 2.2 ;
      RECT 702.96 -35.52 703.28 -31.12 ;
      RECT 702.98 -35.545 703.26 -31.12 ;
      RECT 702.3 -21.24 702.58 2.225 ;
      RECT 702.28 -21.24 702.6 2.2 ;
      RECT 701.6 -35.52 701.92 2.2 ;
      RECT 701.62 -35.545 701.9 2.2 ;
      RECT 700.94 -35.52 701.22 2.225 ;
      RECT 700.92 -35.52 701.24 2.2 ;
      RECT 700.24 -35.52 700.56 2.2 ;
      RECT 700.26 -35.545 700.54 2.2 ;
      RECT 699.58 -35.52 699.86 2.225 ;
      RECT 699.56 -35.52 699.88 2.2 ;
      RECT 698.88 -35.52 699.2 2.2 ;
      RECT 698.9 -35.545 699.18 2.2 ;
      RECT 698.22 -35.52 698.5 2.225 ;
      RECT 698.2 -35.52 698.52 2.2 ;
      RECT 697.52 -35.52 697.84 2.2 ;
      RECT 697.54 -35.545 697.82 2.2 ;
      RECT 696.86 -35.52 697.14 2.225 ;
      RECT 696.84 -35.52 697.16 2.2 ;
      RECT 695.5 -20.56 695.78 2.225 ;
      RECT 695.48 -20.56 695.8 2.2 ;
      RECT 695.44 -35.475 695.76 -30.11 ;
      RECT 695.46 -35.495 695.74 -30.11 ;
      RECT 694.14 -21.24 694.42 2.225 ;
      RECT 694.12 -21.24 694.44 2.2 ;
      RECT 692.78 -25.32 693.06 2.225 ;
      RECT 692.76 -25.32 693.08 2.2 ;
      RECT 691.42 -17.16 691.7 2.225 ;
      RECT 691.4 -17.16 691.72 2.2 ;
      RECT 690.06 -18.52 690.34 2.225 ;
      RECT 690.04 -18.52 690.36 2.2 ;
      RECT 688.7 -18.52 688.98 2.225 ;
      RECT 688.68 -18.52 689 2.2 ;
      RECT 688 -35.52 688.32 -31.12 ;
      RECT 688.02 -35.545 688.3 -31.12 ;
      RECT 687.34 -21.24 687.62 2.225 ;
      RECT 687.32 -21.24 687.64 2.2 ;
      RECT 686.64 -35.52 686.96 2.2 ;
      RECT 686.66 -35.545 686.94 2.2 ;
      RECT 685.98 -35.52 686.26 2.225 ;
      RECT 685.96 -35.52 686.28 2.2 ;
      RECT 685.28 -35.52 685.6 2.2 ;
      RECT 685.3 -35.545 685.58 2.2 ;
      RECT 684.62 -35.52 684.9 2.225 ;
      RECT 684.6 -35.52 684.92 2.2 ;
      RECT 683.92 -35.52 684.24 2.2 ;
      RECT 683.94 -35.545 684.22 2.2 ;
      RECT 683.26 -35.52 683.54 2.225 ;
      RECT 683.24 -35.52 683.56 2.2 ;
      RECT 682.56 -35.52 682.88 2.2 ;
      RECT 682.58 -35.545 682.86 2.2 ;
      RECT 681.9 -35.52 682.18 2.225 ;
      RECT 681.88 -35.52 682.2 2.2 ;
      RECT 680.54 -35.475 680.86 -30.11 ;
      RECT 680.56 -35.495 680.84 -30.11 ;
      RECT 680.54 -20.56 680.82 2.225 ;
      RECT 680.52 -20.56 680.84 2.2 ;
      RECT 679.18 -35.52 679.46 2.225 ;
      RECT 679.16 -35.52 679.48 2.2 ;
      RECT 677.82 -25.32 678.1 2.225 ;
      RECT 677.8 -25.32 678.12 2.2 ;
      RECT 676.46 -17.16 676.74 2.225 ;
      RECT 676.44 -17.16 676.76 2.2 ;
      RECT 675.1 -18.52 675.38 2.225 ;
      RECT 675.08 -18.52 675.4 2.2 ;
      RECT 673.74 -18.52 674.02 2.225 ;
      RECT 673.72 -18.52 674.04 2.2 ;
      RECT 673.04 -35.52 673.36 -31.12 ;
      RECT 673.06 -35.545 673.34 -31.12 ;
      RECT 672.38 -21.24 672.66 2.225 ;
      RECT 672.36 -21.24 672.68 2.2 ;
      RECT 671.68 -35.52 672 2.2 ;
      RECT 671.7 -35.545 671.98 2.2 ;
      RECT 671.02 -35.52 671.3 2.225 ;
      RECT 671 -35.52 671.32 2.2 ;
      RECT 670.32 -35.52 670.64 2.2 ;
      RECT 670.34 -35.545 670.62 2.2 ;
      RECT 669.66 -35.52 669.94 2.225 ;
      RECT 669.64 -35.52 669.96 2.2 ;
      RECT 668.96 -35.52 669.28 2.2 ;
      RECT 668.98 -35.545 669.26 2.2 ;
      RECT 668.3 -35.52 668.58 2.225 ;
      RECT 668.28 -35.52 668.6 2.2 ;
      RECT 667.6 -35.52 667.92 2.2 ;
      RECT 667.62 -35.545 667.9 2.2 ;
      RECT 666.94 -24.64 667.22 2.225 ;
      RECT 666.92 -24.64 667.24 2.2 ;
      RECT 665.64 -35.475 665.96 -30.11 ;
      RECT 665.66 -35.495 665.94 -30.11 ;
      RECT 665.58 -20.56 665.86 2.225 ;
      RECT 665.56 -20.56 665.88 2.2 ;
      RECT 664.22 -35.52 664.5 2.225 ;
      RECT 664.2 -35.52 664.52 2.2 ;
      RECT 662.86 -25.32 663.14 2.225 ;
      RECT 662.84 -25.32 663.16 2.2 ;
      RECT 661.5 -17.16 661.78 2.225 ;
      RECT 661.48 -17.16 661.8 2.2 ;
      RECT 660.14 -18.52 660.42 2.225 ;
      RECT 660.12 -18.52 660.44 2.2 ;
      RECT 658.78 -18.52 659.06 2.225 ;
      RECT 658.76 -18.52 659.08 2.2 ;
      RECT 658.08 -35.52 658.4 -31.12 ;
      RECT 658.1 -35.545 658.38 -31.12 ;
      RECT 657.42 -21.24 657.7 2.225 ;
      RECT 657.4 -21.24 657.72 2.2 ;
      RECT 656.72 -35.52 657.04 2.2 ;
      RECT 656.74 -35.545 657.02 2.2 ;
      RECT 656.06 -35.52 656.34 2.225 ;
      RECT 656.04 -35.52 656.36 2.2 ;
      RECT 655.36 -35.52 655.68 2.2 ;
      RECT 655.38 -35.545 655.66 2.2 ;
      RECT 654.7 -35.52 654.98 2.225 ;
      RECT 654.68 -35.52 655 2.2 ;
      RECT 654 -35.52 654.32 2.2 ;
      RECT 654.02 -35.545 654.3 2.2 ;
      RECT 653.34 -35.52 653.62 2.225 ;
      RECT 653.32 -35.52 653.64 2.2 ;
      RECT 652.64 -35.52 652.96 2.2 ;
      RECT 652.66 -35.545 652.94 2.2 ;
      RECT 651.98 -24.64 652.26 2.225 ;
      RECT 651.96 -24.64 652.28 2.2 ;
      RECT 650.74 -35.475 651.06 -30.11 ;
      RECT 650.76 -35.495 651.04 -30.11 ;
      RECT 650.62 -20.56 650.9 2.225 ;
      RECT 650.6 -20.56 650.92 2.2 ;
      RECT 649.26 -35.52 649.54 2.225 ;
      RECT 649.24 -35.52 649.56 2.2 ;
      RECT 647.9 -25.32 648.18 2.225 ;
      RECT 647.88 -25.32 648.2 2.2 ;
      RECT 646.54 -17.16 646.82 2.225 ;
      RECT 646.52 -17.16 646.84 2.2 ;
      RECT 645.18 -18.52 645.46 2.225 ;
      RECT 645.16 -18.52 645.48 2.2 ;
      RECT 643.82 -18.52 644.1 2.225 ;
      RECT 643.8 -18.52 644.12 2.2 ;
      RECT 643.12 -35.52 643.44 -31.12 ;
      RECT 643.14 -35.545 643.42 -31.12 ;
      RECT 642.46 -21.24 642.74 2.225 ;
      RECT 642.44 -21.24 642.76 2.2 ;
      RECT 641.76 -35.52 642.08 2.2 ;
      RECT 641.78 -35.545 642.06 2.2 ;
      RECT 641.1 -35.52 641.38 2.225 ;
      RECT 641.08 -35.52 641.4 2.2 ;
      RECT 640.4 -35.52 640.72 2.2 ;
      RECT 640.42 -35.545 640.7 2.2 ;
      RECT 639.74 -35.52 640.02 2.225 ;
      RECT 639.72 -35.52 640.04 2.2 ;
      RECT 639.04 -35.52 639.36 2.2 ;
      RECT 639.06 -35.545 639.34 2.2 ;
      RECT 638.38 -35.52 638.66 2.225 ;
      RECT 638.36 -35.52 638.68 2.2 ;
      RECT 637.68 -35.52 638 2.2 ;
      RECT 637.7 -35.545 637.98 2.2 ;
      RECT 637.02 -24.64 637.3 2.225 ;
      RECT 637 -24.64 637.32 2.2 ;
      RECT 635.84 -35.475 636.16 -30.11 ;
      RECT 635.86 -35.495 636.14 -30.11 ;
      RECT 635.66 -20.56 635.94 2.225 ;
      RECT 635.64 -20.56 635.96 2.2 ;
      RECT 634.3 -35.52 634.58 2.225 ;
      RECT 634.28 -35.52 634.6 2.2 ;
      RECT 632.94 -25.32 633.22 2.225 ;
      RECT 632.92 -25.32 633.24 2.2 ;
      RECT 631.58 -17.16 631.86 2.225 ;
      RECT 631.56 -17.16 631.88 2.2 ;
      RECT 630.22 -18.52 630.5 2.225 ;
      RECT 630.2 -18.52 630.52 2.2 ;
      RECT 628.86 -18.52 629.14 2.225 ;
      RECT 628.84 -18.52 629.16 2.2 ;
      RECT 628.16 -35.52 628.48 -31.12 ;
      RECT 628.18 -35.545 628.46 -31.12 ;
      RECT 627.5 -35.52 627.78 2.225 ;
      RECT 627.48 -35.52 627.8 2.2 ;
      RECT 626.8 -35.52 627.12 2.2 ;
      RECT 626.82 -35.545 627.1 2.2 ;
      RECT 626.14 -35.52 626.42 2.225 ;
      RECT 626.12 -35.52 626.44 2.2 ;
      RECT 625.44 -35.52 625.76 2.2 ;
      RECT 625.46 -35.545 625.74 2.2 ;
      RECT 624.78 -35.52 625.06 2.225 ;
      RECT 624.76 -35.52 625.08 2.2 ;
      RECT 624.08 -35.52 624.4 2.2 ;
      RECT 624.1 -35.545 624.38 2.2 ;
      RECT 623.42 -35.52 623.7 2.225 ;
      RECT 623.4 -35.52 623.72 2.2 ;
      RECT 622.72 -35.52 623.04 2.2 ;
      RECT 622.74 -35.545 623.02 2.2 ;
      RECT 622.06 -24.64 622.34 2.225 ;
      RECT 622.04 -24.64 622.36 2.2 ;
      RECT 620.94 -35.475 621.26 -30.11 ;
      RECT 620.96 -35.495 621.24 -30.11 ;
      RECT 620.7 -20.56 620.98 2.225 ;
      RECT 620.68 -20.56 621 2.2 ;
      RECT 619.34 -35.52 619.62 2.225 ;
      RECT 619.32 -35.52 619.64 2.2 ;
      RECT 617.98 -25.32 618.26 2.225 ;
      RECT 617.96 -25.32 618.28 2.2 ;
      RECT 616.62 -17.16 616.9 2.225 ;
      RECT 616.6 -17.16 616.92 2.2 ;
      RECT 615.26 -18.52 615.54 2.225 ;
      RECT 615.24 -18.52 615.56 2.2 ;
      RECT 613.9 -18.52 614.18 2.225 ;
      RECT 613.88 -18.52 614.2 2.2 ;
      RECT 613.2 -35.52 613.52 -31.12 ;
      RECT 613.22 -35.545 613.5 -31.12 ;
      RECT 612.54 -35.52 612.82 2.225 ;
      RECT 612.52 -35.52 612.84 2.2 ;
      RECT 611.84 -35.52 612.16 2.2 ;
      RECT 611.86 -35.545 612.14 2.2 ;
      RECT 611.18 -35.52 611.46 2.225 ;
      RECT 611.16 -35.52 611.48 2.2 ;
      RECT 610.48 -35.52 610.8 2.2 ;
      RECT 610.5 -35.545 610.78 2.2 ;
      RECT 609.82 -35.52 610.1 2.225 ;
      RECT 609.8 -35.52 610.12 2.2 ;
      RECT 609.12 -35.52 609.44 2.2 ;
      RECT 609.14 -35.545 609.42 2.2 ;
      RECT 608.46 -35.52 608.74 2.225 ;
      RECT 608.44 -35.52 608.76 2.2 ;
      RECT 607.76 -35.52 608.08 2.2 ;
      RECT 607.78 -35.545 608.06 2.2 ;
      RECT 607.1 -24.64 607.38 2.225 ;
      RECT 607.08 -24.64 607.4 2.2 ;
      RECT 606.04 -35.475 606.36 -30.11 ;
      RECT 606.06 -35.495 606.34 -30.11 ;
      RECT 605.74 -20.56 606.02 2.225 ;
      RECT 605.72 -20.56 606.04 2.2 ;
      RECT 604.38 -35.52 604.66 2.225 ;
      RECT 604.36 -35.52 604.68 2.2 ;
      RECT 603.02 -25.32 603.3 2.225 ;
      RECT 603 -25.32 603.32 2.2 ;
      RECT 601.66 -17.16 601.94 2.225 ;
      RECT 601.64 -17.16 601.96 2.2 ;
      RECT 600.3 -21.92 600.58 2.225 ;
      RECT 600.28 -21.92 600.6 2.2 ;
      RECT 598.94 -18.52 599.22 2.225 ;
      RECT 598.92 -18.52 599.24 2.2 ;
      RECT 598.24 -35.52 598.56 -31.12 ;
      RECT 598.26 -35.545 598.54 -31.12 ;
      RECT 597.58 -35.52 597.86 2.225 ;
      RECT 597.56 -35.52 597.88 2.2 ;
      RECT 596.88 -35.52 597.2 2.2 ;
      RECT 596.9 -35.545 597.18 2.2 ;
      RECT 596.22 -35.52 596.5 2.225 ;
      RECT 596.2 -35.52 596.52 2.2 ;
      RECT 595.52 -35.52 595.84 2.2 ;
      RECT 595.54 -35.545 595.82 2.2 ;
      RECT 594.86 -35.52 595.14 2.225 ;
      RECT 594.84 -35.52 595.16 2.2 ;
      RECT 594.16 -35.52 594.48 2.2 ;
      RECT 594.18 -35.545 594.46 2.2 ;
      RECT 593.5 -35.52 593.78 2.225 ;
      RECT 593.48 -35.52 593.8 2.2 ;
      RECT 592.8 -35.52 593.12 2.2 ;
      RECT 592.82 -35.545 593.1 2.2 ;
      RECT 592.14 -24.64 592.42 2.225 ;
      RECT 592.12 -24.64 592.44 2.2 ;
      RECT 591.14 -35.475 591.46 -30.11 ;
      RECT 591.16 -35.495 591.44 -30.11 ;
      RECT 590.78 -20.56 591.06 2.225 ;
      RECT 590.76 -20.56 591.08 2.2 ;
      RECT 589.42 -35.52 589.7 2.225 ;
      RECT 589.4 -35.52 589.72 2.2 ;
      RECT 588.06 -25.32 588.34 2.225 ;
      RECT 588.04 -25.32 588.36 2.2 ;
      RECT 586.7 -17.84 586.98 2.225 ;
      RECT 586.68 -17.84 587 2.2 ;
      RECT 585.34 -21.92 585.62 2.225 ;
      RECT 585.32 -21.92 585.64 2.2 ;
      RECT 583.98 -18.52 584.26 2.225 ;
      RECT 583.96 -18.52 584.28 2.2 ;
      RECT 583.28 -35.52 583.6 -31.12 ;
      RECT 583.3 -35.545 583.58 -31.12 ;
      RECT 582.62 -35.52 582.9 2.225 ;
      RECT 582.6 -35.52 582.92 2.2 ;
      RECT 581.92 -35.52 582.24 2.2 ;
      RECT 581.94 -35.545 582.22 2.2 ;
      RECT 581.26 -35.52 581.54 2.225 ;
      RECT 581.24 -35.52 581.56 2.2 ;
      RECT 580.56 -35.52 580.88 2.2 ;
      RECT 580.58 -35.545 580.86 2.2 ;
      RECT 579.9 -35.52 580.18 2.225 ;
      RECT 579.88 -35.52 580.2 2.2 ;
      RECT 579.2 -35.52 579.52 2.2 ;
      RECT 579.22 -35.545 579.5 2.2 ;
      RECT 578.54 -35.52 578.82 2.225 ;
      RECT 578.52 -35.52 578.84 2.2 ;
      RECT 577.84 -35.52 578.16 2.2 ;
      RECT 577.86 -35.545 578.14 2.2 ;
      RECT 577.18 -24.64 577.46 2.225 ;
      RECT 577.16 -24.64 577.48 2.2 ;
      RECT 576.24 -35.475 576.56 -30.11 ;
      RECT 576.26 -35.495 576.54 -30.11 ;
      RECT 575.82 -20.56 576.1 2.225 ;
      RECT 575.8 -20.56 576.12 2.2 ;
      RECT 574.46 -35.52 574.74 2.225 ;
      RECT 574.44 -35.52 574.76 2.2 ;
      RECT 573.1 -17.16 573.38 2.225 ;
      RECT 573.08 -17.16 573.4 2.2 ;
      RECT 571.74 -17.84 572.02 2.225 ;
      RECT 571.72 -17.84 572.04 2.2 ;
      RECT 570.38 -21.92 570.66 2.225 ;
      RECT 570.36 -21.92 570.68 2.2 ;
      RECT 569.02 -18.52 569.3 2.225 ;
      RECT 569 -18.52 569.32 2.2 ;
      RECT 568.32 -35.52 568.64 -31.12 ;
      RECT 568.34 -35.545 568.62 -31.12 ;
      RECT 567.66 -35.52 567.94 2.225 ;
      RECT 567.64 -35.52 567.96 2.2 ;
      RECT 566.96 -35.52 567.28 2.2 ;
      RECT 566.98 -35.545 567.26 2.2 ;
      RECT 566.3 -35.52 566.58 2.225 ;
      RECT 566.28 -35.52 566.6 2.2 ;
      RECT 565.6 -35.52 565.92 2.2 ;
      RECT 565.62 -35.545 565.9 2.2 ;
      RECT 564.94 -35.52 565.22 2.225 ;
      RECT 564.92 -35.52 565.24 2.2 ;
      RECT 564.24 -35.52 564.56 2.2 ;
      RECT 564.26 -35.545 564.54 2.2 ;
      RECT 563.58 -35.52 563.86 2.225 ;
      RECT 563.56 -35.52 563.88 2.2 ;
      RECT 562.88 -35.52 563.2 2.2 ;
      RECT 562.9 -35.545 563.18 2.2 ;
      RECT 562.22 -24.64 562.5 2.225 ;
      RECT 562.2 -24.64 562.52 2.2 ;
      RECT 561.34 -35.475 561.66 -30.11 ;
      RECT 561.36 -35.495 561.64 -30.11 ;
      RECT 560.86 -20.56 561.14 2.225 ;
      RECT 560.84 -20.56 561.16 2.2 ;
      RECT 559.5 -25.32 559.78 2.225 ;
      RECT 559.48 -25.32 559.8 2.2 ;
      RECT 558.14 -17.16 558.42 2.225 ;
      RECT 558.12 -17.16 558.44 2.2 ;
      RECT 556.78 -17.84 557.06 2.225 ;
      RECT 556.76 -17.84 557.08 2.2 ;
      RECT 555.42 -21.92 555.7 2.225 ;
      RECT 555.4 -21.92 555.72 2.2 ;
      RECT 554.06 -18.52 554.34 2.225 ;
      RECT 554.04 -18.52 554.36 2.2 ;
      RECT 553.36 -35.52 553.68 -31.12 ;
      RECT 553.38 -35.545 553.66 -31.12 ;
      RECT 552.7 -35.52 552.98 2.225 ;
      RECT 552.68 -35.52 553 2.2 ;
      RECT 552 -35.52 552.32 2.2 ;
      RECT 552.02 -35.545 552.3 2.2 ;
      RECT 551.34 -35.52 551.62 2.225 ;
      RECT 551.32 -35.52 551.64 2.2 ;
      RECT 550.64 -35.52 550.96 2.2 ;
      RECT 550.66 -35.545 550.94 2.2 ;
      RECT 549.98 -35.52 550.26 2.225 ;
      RECT 549.96 -35.52 550.28 2.2 ;
      RECT 549.28 -35.52 549.6 2.2 ;
      RECT 549.3 -35.545 549.58 2.2 ;
      RECT 548.62 -35.52 548.9 2.225 ;
      RECT 548.6 -35.52 548.92 2.2 ;
      RECT 547.92 -35.52 548.24 2.2 ;
      RECT 547.94 -35.545 548.22 2.2 ;
      RECT 547.26 -24.64 547.54 2.225 ;
      RECT 547.24 -24.64 547.56 2.2 ;
      RECT 546.44 -35.475 546.76 -30.11 ;
      RECT 546.46 -35.495 546.74 -30.11 ;
      RECT 545.9 -20.56 546.18 2.225 ;
      RECT 545.88 -20.56 546.2 2.2 ;
      RECT 544.54 -25.32 544.82 2.225 ;
      RECT 544.52 -25.32 544.84 2.2 ;
      RECT 543.18 -17.16 543.46 2.225 ;
      RECT 543.16 -17.16 543.48 2.2 ;
      RECT 541.82 -17.84 542.1 2.225 ;
      RECT 541.8 -17.84 542.12 2.2 ;
      RECT 540.46 -21.92 540.74 2.225 ;
      RECT 540.44 -21.92 540.76 2.2 ;
      RECT 539.1 -18.52 539.38 2.225 ;
      RECT 539.08 -18.52 539.4 2.2 ;
      RECT 538.4 -35.52 538.72 -31.12 ;
      RECT 538.42 -35.545 538.7 -31.12 ;
      RECT 537.74 -35.52 538.02 2.225 ;
      RECT 537.72 -35.52 538.04 2.2 ;
      RECT 537.04 -35.52 537.36 2.2 ;
      RECT 537.06 -35.545 537.34 2.2 ;
      RECT 536.38 -35.52 536.66 2.225 ;
      RECT 536.36 -35.52 536.68 2.2 ;
      RECT 535.68 -35.52 536 2.2 ;
      RECT 535.7 -35.545 535.98 2.2 ;
      RECT 535.02 -35.52 535.3 2.225 ;
      RECT 535 -35.52 535.32 2.2 ;
      RECT 534.32 -35.52 534.64 2.2 ;
      RECT 534.34 -35.545 534.62 2.2 ;
      RECT 533.66 -35.52 533.94 2.225 ;
      RECT 533.64 -35.52 533.96 2.2 ;
      RECT 532.96 -35.52 533.28 2.2 ;
      RECT 532.98 -35.545 533.26 2.2 ;
      RECT 532.3 -24.64 532.58 2.225 ;
      RECT 532.28 -24.64 532.6 2.2 ;
      RECT 531.54 -35.475 531.86 -30.11 ;
      RECT 531.56 -35.495 531.84 -30.11 ;
      RECT 530.94 -20.56 531.22 2.225 ;
      RECT 530.92 -20.56 531.24 2.2 ;
      RECT 529.58 -25.32 529.86 2.225 ;
      RECT 529.56 -25.32 529.88 2.2 ;
      RECT 528.22 -17.16 528.5 2.225 ;
      RECT 528.2 -17.16 528.52 2.2 ;
      RECT 526.86 -17.84 527.14 2.225 ;
      RECT 526.84 -17.84 527.16 2.2 ;
      RECT 525.5 -21.92 525.78 2.225 ;
      RECT 525.48 -21.92 525.8 2.2 ;
      RECT 524.14 -18.52 524.42 2.225 ;
      RECT 524.12 -18.52 524.44 2.2 ;
      RECT 523.44 -35.52 523.76 -31.12 ;
      RECT 523.46 -35.545 523.74 -31.12 ;
      RECT 522.78 -35.52 523.06 2.225 ;
      RECT 522.76 -35.52 523.08 2.2 ;
      RECT 522.08 -35.52 522.4 2.2 ;
      RECT 522.1 -35.545 522.38 2.2 ;
      RECT 521.42 -35.52 521.7 2.225 ;
      RECT 521.4 -35.52 521.72 2.2 ;
      RECT 520.72 -35.52 521.04 2.2 ;
      RECT 520.74 -35.545 521.02 2.2 ;
      RECT 520.06 -35.52 520.34 2.225 ;
      RECT 520.04 -35.52 520.36 2.2 ;
      RECT 519.36 -35.52 519.68 2.2 ;
      RECT 519.38 -35.545 519.66 2.2 ;
      RECT 518.7 -35.52 518.98 2.225 ;
      RECT 518.68 -35.52 519 2.2 ;
      RECT 518 -35.52 518.32 2.2 ;
      RECT 518.02 -35.545 518.3 2.2 ;
      RECT 517.34 -24.64 517.62 2.225 ;
      RECT 517.32 -24.64 517.64 2.2 ;
      RECT 516.64 -35.475 516.96 -30.11 ;
      RECT 516.66 -35.495 516.94 -30.11 ;
      RECT 515.98 -21.24 516.26 2.225 ;
      RECT 515.96 -21.24 516.28 2.2 ;
      RECT 514.62 -25.32 514.9 2.225 ;
      RECT 514.6 -25.32 514.92 2.2 ;
      RECT 513.26 -17.16 513.54 2.225 ;
      RECT 513.24 -17.16 513.56 2.2 ;
      RECT 511.9 -17.84 512.18 2.225 ;
      RECT 511.88 -17.84 512.2 2.2 ;
      RECT 510.54 -21.92 510.82 2.225 ;
      RECT 510.52 -21.92 510.84 2.2 ;
      RECT 509.18 -18.52 509.46 2.225 ;
      RECT 509.16 -18.52 509.48 2.2 ;
      RECT 508.48 -35.52 508.8 -31.12 ;
      RECT 508.5 -35.545 508.78 -31.12 ;
      RECT 507.82 -35.52 508.1 2.225 ;
      RECT 507.8 -35.52 508.12 2.2 ;
      RECT 507.12 -35.52 507.44 2.2 ;
      RECT 507.14 -35.545 507.42 2.2 ;
      RECT 506.46 -35.52 506.74 2.225 ;
      RECT 506.44 -35.52 506.76 2.2 ;
      RECT 505.76 -35.52 506.08 2.2 ;
      RECT 505.78 -35.545 506.06 2.2 ;
      RECT 505.1 -35.52 505.38 2.225 ;
      RECT 505.08 -35.52 505.4 2.2 ;
      RECT 504.4 -35.52 504.72 2.2 ;
      RECT 504.42 -35.545 504.7 2.2 ;
      RECT 503.74 -35.52 504.02 2.225 ;
      RECT 503.72 -35.52 504.04 2.2 ;
      RECT 502.38 -20.56 502.66 2.225 ;
      RECT 502.36 -20.56 502.68 2.2 ;
      RECT 501.74 -35.475 502.06 -30.11 ;
      RECT 501.76 -35.495 502.04 -30.11 ;
      RECT 501.02 -21.24 501.3 2.225 ;
      RECT 501 -21.24 501.32 2.2 ;
      RECT 499.66 -25.32 499.94 2.225 ;
      RECT 499.64 -25.32 499.96 2.2 ;
      RECT 498.3 -17.16 498.58 2.225 ;
      RECT 498.28 -17.16 498.6 2.2 ;
      RECT 496.94 -17.84 497.22 2.225 ;
      RECT 496.92 -17.84 497.24 2.2 ;
      RECT 495.58 -21.92 495.86 2.225 ;
      RECT 495.56 -21.92 495.88 2.2 ;
      RECT 494.22 -18.52 494.5 2.225 ;
      RECT 494.2 -18.52 494.52 2.2 ;
      RECT 493.52 -35.52 493.84 -31.12 ;
      RECT 493.54 -35.545 493.82 -31.12 ;
      RECT 492.86 -35.52 493.14 2.225 ;
      RECT 492.84 -35.52 493.16 2.2 ;
      RECT 492.16 -35.52 492.48 2.2 ;
      RECT 492.18 -35.545 492.46 2.2 ;
      RECT 491.5 -35.52 491.78 2.225 ;
      RECT 491.48 -35.52 491.8 2.2 ;
      RECT 490.8 -35.52 491.12 2.2 ;
      RECT 490.82 -35.545 491.1 2.2 ;
      RECT 490.14 -35.52 490.42 2.225 ;
      RECT 490.12 -35.52 490.44 2.2 ;
      RECT 489.44 -35.52 489.76 2.2 ;
      RECT 489.46 -35.545 489.74 2.2 ;
      RECT 488.78 -35.52 489.06 2.225 ;
      RECT 488.76 -35.52 489.08 2.2 ;
      RECT 487.42 -20.56 487.7 2.225 ;
      RECT 487.4 -20.56 487.72 2.2 ;
      RECT 486.84 -35.475 487.16 -30.11 ;
      RECT 486.86 -35.495 487.14 -30.11 ;
      RECT 486.06 -21.24 486.34 2.225 ;
      RECT 486.04 -21.24 486.36 2.2 ;
      RECT 484.7 -25.32 484.98 2.225 ;
      RECT 484.68 -25.32 485 2.2 ;
      RECT 483.34 -17.16 483.62 2.225 ;
      RECT 483.32 -17.16 483.64 2.2 ;
      RECT 481.98 -17.84 482.26 2.225 ;
      RECT 481.96 -17.84 482.28 2.2 ;
      RECT 480.62 -21.92 480.9 2.225 ;
      RECT 480.6 -21.92 480.92 2.2 ;
      RECT 479.26 -18.52 479.54 2.225 ;
      RECT 479.24 -18.52 479.56 2.2 ;
      RECT 478.56 -35.52 478.88 -31.12 ;
      RECT 478.58 -35.545 478.86 -31.12 ;
      RECT 477.9 -35.52 478.18 2.225 ;
      RECT 477.88 -35.52 478.2 2.2 ;
      RECT 477.2 -35.52 477.52 2.2 ;
      RECT 477.22 -35.545 477.5 2.2 ;
      RECT 476.54 -35.52 476.82 2.225 ;
      RECT 476.52 -35.52 476.84 2.2 ;
      RECT 475.84 -35.52 476.16 2.2 ;
      RECT 475.86 -35.545 476.14 2.2 ;
      RECT 475.18 -35.52 475.46 2.225 ;
      RECT 475.16 -35.52 475.48 2.2 ;
      RECT 474.48 -35.52 474.8 2.2 ;
      RECT 474.5 -35.545 474.78 2.2 ;
      RECT 473.82 -35.52 474.1 2.225 ;
      RECT 473.8 -35.52 474.12 2.2 ;
      RECT 472.46 -20.56 472.74 2.225 ;
      RECT 472.44 -20.56 472.76 2.2 ;
      RECT 471.94 -35.475 472.26 -30.11 ;
      RECT 471.96 -35.495 472.24 -30.11 ;
      RECT 471.1 -21.24 471.38 2.225 ;
      RECT 471.08 -21.24 471.4 2.2 ;
      RECT 469.74 -25.32 470.02 2.225 ;
      RECT 469.72 -25.32 470.04 2.2 ;
      RECT 468.38 -17.16 468.66 2.225 ;
      RECT 468.36 -17.16 468.68 2.2 ;
      RECT 467.02 -17.84 467.3 2.225 ;
      RECT 467 -17.84 467.32 2.2 ;
      RECT 465.66 -18.52 465.94 2.225 ;
      RECT 465.64 -18.52 465.96 2.2 ;
      RECT 464.3 -21.24 464.58 2.225 ;
      RECT 464.28 -21.24 464.6 2.2 ;
      RECT 463.6 -35.52 463.92 2.2 ;
      RECT 463.62 -35.545 463.9 2.2 ;
      RECT 462.94 -35.52 463.22 2.225 ;
      RECT 462.92 -35.52 463.24 2.2 ;
      RECT 462.24 -35.52 462.56 2.2 ;
      RECT 462.26 -35.545 462.54 2.2 ;
      RECT 461.58 -35.52 461.86 2.225 ;
      RECT 461.56 -35.52 461.88 2.2 ;
      RECT 460.88 -35.52 461.2 2.2 ;
      RECT 460.9 -35.545 461.18 2.2 ;
      RECT 460.22 -35.52 460.5 2.225 ;
      RECT 460.2 -35.52 460.52 2.2 ;
      RECT 459.52 -35.52 459.84 2.2 ;
      RECT 459.54 -35.545 459.82 2.2 ;
      RECT 458.86 -35.52 459.14 2.225 ;
      RECT 458.84 -35.52 459.16 2.2 ;
      RECT 457.5 -20.56 457.78 2.225 ;
      RECT 457.48 -20.56 457.8 2.2 ;
      RECT 457.04 -35.475 457.36 -30.11 ;
      RECT 457.06 -35.495 457.34 -30.11 ;
      RECT 456.14 -21.24 456.42 2.225 ;
      RECT 456.12 -21.24 456.44 2.2 ;
      RECT 454.78 -25.32 455.06 2.225 ;
      RECT 454.76 -25.32 455.08 2.2 ;
      RECT 453.42 -17.16 453.7 2.225 ;
      RECT 453.4 -17.16 453.72 2.2 ;
      RECT 452.06 -17.84 452.34 2.225 ;
      RECT 452.04 -17.84 452.36 2.2 ;
      RECT 450.7 -18.52 450.98 2.225 ;
      RECT 450.68 -18.52 451 2.2 ;
      RECT 450 -35.52 450.32 -31.12 ;
      RECT 450.02 -35.545 450.3 -31.12 ;
      RECT 449.34 -21.24 449.62 2.225 ;
      RECT 449.32 -21.24 449.64 2.2 ;
      RECT 448.64 -35.52 448.96 2.2 ;
      RECT 448.66 -35.545 448.94 2.2 ;
      RECT 447.98 -35.52 448.26 2.225 ;
      RECT 447.96 -35.52 448.28 2.2 ;
      RECT 447.28 -35.52 447.6 2.2 ;
      RECT 447.3 -35.545 447.58 2.2 ;
      RECT 446.62 -35.52 446.9 2.225 ;
      RECT 446.6 -35.52 446.92 2.2 ;
      RECT 445.92 -35.52 446.24 2.2 ;
      RECT 445.94 -35.545 446.22 2.2 ;
      RECT 445.26 -35.52 445.54 2.225 ;
      RECT 445.24 -35.52 445.56 2.2 ;
      RECT 444.56 -35.52 444.88 2.2 ;
      RECT 444.58 -35.545 444.86 2.2 ;
      RECT 443.9 -35.52 444.18 2.225 ;
      RECT 443.88 -35.52 444.2 2.2 ;
      RECT 442.54 -20.56 442.82 2.225 ;
      RECT 442.52 -20.56 442.84 2.2 ;
      RECT 442.14 -35.475 442.46 -30.11 ;
      RECT 442.16 -35.495 442.44 -30.11 ;
      RECT 441.18 -21.24 441.46 2.225 ;
      RECT 441.16 -21.24 441.48 2.2 ;
      RECT 439.82 -25.32 440.1 2.225 ;
      RECT 439.8 -25.32 440.12 2.2 ;
      RECT 438.46 -17.16 438.74 2.225 ;
      RECT 438.44 -17.16 438.76 2.2 ;
      RECT 437.1 -17.84 437.38 2.225 ;
      RECT 437.08 -17.84 437.4 2.2 ;
      RECT 435.74 -18.52 436.02 2.225 ;
      RECT 435.72 -18.52 436.04 2.2 ;
      RECT 435.04 -35.52 435.36 -31.12 ;
      RECT 435.06 -35.545 435.34 -31.12 ;
      RECT 434.38 -21.24 434.66 2.225 ;
      RECT 434.36 -21.24 434.68 2.2 ;
      RECT 433.68 -35.52 434 2.2 ;
      RECT 433.7 -35.545 433.98 2.2 ;
      RECT 433.02 -35.52 433.3 2.225 ;
      RECT 433 -35.52 433.32 2.2 ;
      RECT 432.32 -35.52 432.64 2.2 ;
      RECT 432.34 -35.545 432.62 2.2 ;
      RECT 431.66 -35.52 431.94 2.225 ;
      RECT 431.64 -35.52 431.96 2.2 ;
      RECT 430.96 -35.52 431.28 2.2 ;
      RECT 430.98 -35.545 431.26 2.2 ;
      RECT 430.3 -35.52 430.58 2.225 ;
      RECT 430.28 -35.52 430.6 2.2 ;
      RECT 429.6 -35.52 429.92 2.2 ;
      RECT 429.62 -35.545 429.9 2.2 ;
      RECT 428.94 -35.52 429.22 2.225 ;
      RECT 428.92 -35.52 429.24 2.2 ;
      RECT 427.58 -20.56 427.86 2.225 ;
      RECT 427.56 -20.56 427.88 2.2 ;
      RECT 427.24 -35.475 427.56 -30.11 ;
      RECT 427.26 -35.495 427.54 -30.11 ;
      RECT 426.22 -21.24 426.5 2.225 ;
      RECT 426.2 -21.24 426.52 2.2 ;
      RECT 424.86 -25.32 425.14 2.225 ;
      RECT 424.84 -25.32 425.16 2.2 ;
      RECT 423.5 -17.16 423.78 2.225 ;
      RECT 423.48 -17.16 423.8 2.2 ;
      RECT 422.14 -18.52 422.42 2.225 ;
      RECT 422.12 -18.52 422.44 2.2 ;
      RECT 420.78 -18.52 421.06 2.225 ;
      RECT 420.76 -18.52 421.08 2.2 ;
      RECT 420.08 -35.52 420.4 -31.12 ;
      RECT 420.1 -35.545 420.38 -31.12 ;
      RECT 419.42 -21.24 419.7 2.225 ;
      RECT 419.4 -21.24 419.72 2.2 ;
      RECT 418.72 -35.52 419.04 2.2 ;
      RECT 418.74 -35.545 419.02 2.2 ;
      RECT 418.06 -35.52 418.34 2.225 ;
      RECT 418.04 -35.52 418.36 2.2 ;
      RECT 417.36 -35.52 417.68 2.2 ;
      RECT 417.38 -35.545 417.66 2.2 ;
      RECT 416.7 -35.52 416.98 2.225 ;
      RECT 416.68 -35.52 417 2.2 ;
      RECT 416 -35.52 416.32 2.2 ;
      RECT 416.02 -35.545 416.3 2.2 ;
      RECT 415.34 -35.52 415.62 2.225 ;
      RECT 415.32 -35.52 415.64 2.2 ;
      RECT 414.64 -35.52 414.96 2.2 ;
      RECT 414.66 -35.545 414.94 2.2 ;
      RECT 413.98 -35.52 414.26 2.225 ;
      RECT 413.96 -35.52 414.28 2.2 ;
      RECT 412.62 -20.56 412.9 2.225 ;
      RECT 412.6 -20.56 412.92 2.2 ;
      RECT 412.34 -35.475 412.66 -30.11 ;
      RECT 412.36 -35.495 412.64 -30.11 ;
      RECT 411.26 -21.24 411.54 2.225 ;
      RECT 411.24 -21.24 411.56 2.2 ;
      RECT 409.9 -25.32 410.18 2.225 ;
      RECT 409.88 -25.32 410.2 2.2 ;
      RECT 408.54 -17.16 408.82 2.225 ;
      RECT 408.52 -17.16 408.84 2.2 ;
      RECT 407.18 -18.52 407.46 2.225 ;
      RECT 407.16 -18.52 407.48 2.2 ;
      RECT 405.82 -18.52 406.1 2.225 ;
      RECT 405.8 -18.52 406.12 2.2 ;
      RECT 405.12 -35.52 405.44 -31.12 ;
      RECT 405.14 -35.545 405.42 -31.12 ;
      RECT 404.46 -21.24 404.74 2.225 ;
      RECT 404.44 -21.24 404.76 2.2 ;
      RECT 403.76 -35.52 404.08 2.2 ;
      RECT 403.78 -35.545 404.06 2.2 ;
      RECT 403.1 -35.52 403.38 2.225 ;
      RECT 403.08 -35.52 403.4 2.2 ;
      RECT 402.4 -35.52 402.72 2.2 ;
      RECT 402.42 -35.545 402.7 2.2 ;
      RECT 401.74 -35.52 402.02 2.225 ;
      RECT 401.72 -35.52 402.04 2.2 ;
      RECT 401.04 -35.52 401.36 2.2 ;
      RECT 401.06 -35.545 401.34 2.2 ;
      RECT 400.38 -35.52 400.66 2.225 ;
      RECT 400.36 -35.52 400.68 2.2 ;
      RECT 399.68 -35.52 400 2.2 ;
      RECT 399.7 -35.545 399.98 2.2 ;
      RECT 399.02 -35.52 399.3 2.225 ;
      RECT 399 -35.52 399.32 2.2 ;
      RECT 397.66 -20.56 397.94 2.225 ;
      RECT 397.64 -20.56 397.96 2.2 ;
      RECT 397.44 -35.475 397.76 -30.11 ;
      RECT 397.46 -35.495 397.74 -30.11 ;
      RECT 396.3 -21.24 396.58 2.225 ;
      RECT 396.28 -21.24 396.6 2.2 ;
      RECT 394.94 -25.32 395.22 2.225 ;
      RECT 394.92 -25.32 395.24 2.2 ;
      RECT 393.58 -17.16 393.86 2.225 ;
      RECT 393.56 -17.16 393.88 2.2 ;
      RECT 392.22 -18.52 392.5 2.225 ;
      RECT 392.2 -18.52 392.52 2.2 ;
      RECT 390.86 -18.52 391.14 2.225 ;
      RECT 390.84 -18.52 391.16 2.2 ;
      RECT 390.16 -35.52 390.48 -31.12 ;
      RECT 390.18 -35.545 390.46 -31.12 ;
      RECT 389.5 -21.24 389.78 2.225 ;
      RECT 389.48 -21.24 389.8 2.2 ;
      RECT 388.8 -35.52 389.12 2.2 ;
      RECT 388.82 -35.545 389.1 2.2 ;
      RECT 388.14 -35.52 388.42 2.225 ;
      RECT 388.12 -35.52 388.44 2.2 ;
      RECT 387.44 -35.52 387.76 2.2 ;
      RECT 387.46 -35.545 387.74 2.2 ;
      RECT 386.78 -35.52 387.06 2.225 ;
      RECT 386.76 -35.52 387.08 2.2 ;
      RECT 386.08 -35.52 386.4 2.2 ;
      RECT 386.1 -35.545 386.38 2.2 ;
      RECT 385.42 -35.52 385.7 2.225 ;
      RECT 385.4 -35.52 385.72 2.2 ;
      RECT 384.72 -35.52 385.04 2.2 ;
      RECT 384.74 -35.545 385.02 2.2 ;
      RECT 384.06 -35.52 384.34 2.225 ;
      RECT 384.04 -35.52 384.36 2.2 ;
      RECT 382.7 -20.56 382.98 2.225 ;
      RECT 382.68 -20.56 383 2.2 ;
      RECT 382.54 -35.475 382.86 -30.11 ;
      RECT 382.56 -35.495 382.84 -30.11 ;
      RECT 381.34 -21.24 381.62 2.225 ;
      RECT 381.32 -21.24 381.64 2.2 ;
      RECT 379.98 -25.32 380.26 2.225 ;
      RECT 379.96 -25.32 380.28 2.2 ;
      RECT 378.62 -17.16 378.9 2.225 ;
      RECT 378.6 -17.16 378.92 2.2 ;
      RECT 377.26 -18.52 377.54 2.225 ;
      RECT 377.24 -18.52 377.56 2.2 ;
      RECT 375.9 -18.52 376.18 2.225 ;
      RECT 375.88 -18.52 376.2 2.2 ;
      RECT 375.2 -35.52 375.52 -31.12 ;
      RECT 375.22 -35.545 375.5 -31.12 ;
      RECT 374.54 -21.24 374.82 2.225 ;
      RECT 374.52 -21.24 374.84 2.2 ;
      RECT 373.84 -35.52 374.16 2.2 ;
      RECT 373.86 -35.545 374.14 2.2 ;
      RECT 373.18 -35.52 373.46 2.225 ;
      RECT 373.16 -35.52 373.48 2.2 ;
      RECT 372.48 -35.52 372.8 2.2 ;
      RECT 372.5 -35.545 372.78 2.2 ;
      RECT 371.82 -35.52 372.1 2.225 ;
      RECT 371.8 -35.52 372.12 2.2 ;
      RECT 371.12 -35.52 371.44 2.2 ;
      RECT 371.14 -35.545 371.42 2.2 ;
      RECT 370.46 -35.52 370.74 2.225 ;
      RECT 370.44 -35.52 370.76 2.2 ;
      RECT 369.76 -35.52 370.08 2.2 ;
      RECT 369.78 -35.545 370.06 2.2 ;
      RECT 369.1 -35.52 369.38 2.225 ;
      RECT 369.08 -35.52 369.4 2.2 ;
      RECT 367.74 -20.56 368.02 2.225 ;
      RECT 367.72 -20.56 368.04 2.2 ;
      RECT 367.64 -35.475 367.96 -30.11 ;
      RECT 367.66 -35.495 367.94 -30.11 ;
      RECT 366.38 -21.24 366.66 2.225 ;
      RECT 366.36 -21.24 366.68 2.2 ;
      RECT 365.02 -25.32 365.3 2.225 ;
      RECT 365 -25.32 365.32 2.2 ;
      RECT 363.66 -17.16 363.94 2.225 ;
      RECT 363.64 -17.16 363.96 2.2 ;
      RECT 362.3 -18.52 362.58 2.225 ;
      RECT 362.28 -18.52 362.6 2.2 ;
      RECT 360.94 -18.52 361.22 2.225 ;
      RECT 360.92 -18.52 361.24 2.2 ;
      RECT 360.24 -35.52 360.56 -31.12 ;
      RECT 360.26 -35.545 360.54 -31.12 ;
      RECT 359.58 -21.24 359.86 2.225 ;
      RECT 359.56 -21.24 359.88 2.2 ;
      RECT 358.88 -35.52 359.2 2.2 ;
      RECT 358.9 -35.545 359.18 2.2 ;
      RECT 358.22 -35.52 358.5 2.225 ;
      RECT 358.2 -35.52 358.52 2.2 ;
      RECT 357.52 -35.52 357.84 2.2 ;
      RECT 357.54 -35.545 357.82 2.2 ;
      RECT 356.86 -35.52 357.14 2.225 ;
      RECT 356.84 -35.52 357.16 2.2 ;
      RECT 356.16 -35.52 356.48 2.2 ;
      RECT 356.18 -35.545 356.46 2.2 ;
      RECT 355.5 -35.52 355.78 2.225 ;
      RECT 355.48 -35.52 355.8 2.2 ;
      RECT 354.8 -35.52 355.12 2.2 ;
      RECT 354.82 -35.545 355.1 2.2 ;
      RECT 354.14 -35.52 354.42 2.225 ;
      RECT 354.12 -35.52 354.44 2.2 ;
      RECT 352.78 -20.56 353.06 2.225 ;
      RECT 352.76 -20.56 353.08 2.2 ;
      RECT 352.74 -35.475 353.06 -30.11 ;
      RECT 352.76 -35.495 353.04 -30.11 ;
      RECT 351.42 -35.52 351.7 2.225 ;
      RECT 351.4 -35.52 351.72 2.2 ;
      RECT 350.06 -25.32 350.34 2.225 ;
      RECT 350.04 -25.32 350.36 2.2 ;
      RECT 348.7 -17.16 348.98 2.225 ;
      RECT 348.68 -17.16 349 2.2 ;
      RECT 347.34 -18.52 347.62 2.225 ;
      RECT 347.32 -18.52 347.64 2.2 ;
      RECT 345.98 -18.52 346.26 2.225 ;
      RECT 345.96 -18.52 346.28 2.2 ;
      RECT 345.28 -35.52 345.6 -31.12 ;
      RECT 345.3 -35.545 345.58 -31.12 ;
      RECT 344.62 -21.24 344.9 2.225 ;
      RECT 344.6 -21.24 344.92 2.2 ;
      RECT 343.92 -35.52 344.24 2.2 ;
      RECT 343.94 -35.545 344.22 2.2 ;
      RECT 343.26 -35.52 343.54 2.225 ;
      RECT 343.24 -35.52 343.56 2.2 ;
      RECT 342.56 -35.52 342.88 2.2 ;
      RECT 342.58 -35.545 342.86 2.2 ;
      RECT 341.9 -35.52 342.18 2.225 ;
      RECT 341.88 -35.52 342.2 2.2 ;
      RECT 341.2 -35.52 341.52 2.2 ;
      RECT 341.22 -35.545 341.5 2.2 ;
      RECT 340.54 -35.52 340.82 2.225 ;
      RECT 340.52 -35.52 340.84 2.2 ;
      RECT 339.84 -35.52 340.16 2.2 ;
      RECT 339.86 -35.545 340.14 2.2 ;
      RECT 339.18 -35.52 339.46 2.225 ;
      RECT 339.16 -35.52 339.48 2.2 ;
      RECT 337.84 -35.475 338.16 -30.11 ;
      RECT 337.86 -35.495 338.14 -30.11 ;
      RECT 337.82 -20.56 338.1 2.225 ;
      RECT 337.8 -20.56 338.12 2.2 ;
      RECT 336.46 -35.52 336.74 2.225 ;
      RECT 336.44 -35.52 336.76 2.2 ;
      RECT 335.1 -25.32 335.38 2.225 ;
      RECT 335.08 -25.32 335.4 2.2 ;
      RECT 333.74 -17.16 334.02 2.225 ;
      RECT 333.72 -17.16 334.04 2.2 ;
      RECT 332.38 -18.52 332.66 2.225 ;
      RECT 332.36 -18.52 332.68 2.2 ;
      RECT 331.02 -18.52 331.3 2.225 ;
      RECT 331 -18.52 331.32 2.2 ;
      RECT 330.32 -35.52 330.64 -31.12 ;
      RECT 330.34 -35.545 330.62 -31.12 ;
      RECT 329.66 -21.24 329.94 2.225 ;
      RECT 329.64 -21.24 329.96 2.2 ;
      RECT 328.96 -35.52 329.28 2.2 ;
      RECT 328.98 -35.545 329.26 2.2 ;
      RECT 328.3 -35.52 328.58 2.225 ;
      RECT 328.28 -35.52 328.6 2.2 ;
      RECT 327.6 -35.52 327.92 2.2 ;
      RECT 327.62 -35.545 327.9 2.2 ;
      RECT 326.94 -35.52 327.22 2.225 ;
      RECT 326.92 -35.52 327.24 2.2 ;
      RECT 326.24 -35.52 326.56 2.2 ;
      RECT 326.26 -35.545 326.54 2.2 ;
      RECT 325.58 -35.52 325.86 2.225 ;
      RECT 325.56 -35.52 325.88 2.2 ;
      RECT 324.88 -35.52 325.2 2.2 ;
      RECT 324.9 -35.545 325.18 2.2 ;
      RECT 324.22 -24.64 324.5 2.225 ;
      RECT 324.2 -24.64 324.52 2.2 ;
      RECT 322.94 -35.475 323.26 -30.11 ;
      RECT 322.96 -35.495 323.24 -30.11 ;
      RECT 322.86 -20.56 323.14 2.225 ;
      RECT 322.84 -20.56 323.16 2.2 ;
      RECT 321.5 -35.52 321.78 2.225 ;
      RECT 321.48 -35.52 321.8 2.2 ;
      RECT 320.14 -25.32 320.42 2.225 ;
      RECT 320.12 -25.32 320.44 2.2 ;
      RECT 318.78 -17.16 319.06 2.225 ;
      RECT 318.76 -17.16 319.08 2.2 ;
      RECT 317.42 -18.52 317.7 2.225 ;
      RECT 317.4 -18.52 317.72 2.2 ;
      RECT 316.06 -18.52 316.34 2.225 ;
      RECT 316.04 -18.52 316.36 2.2 ;
      RECT 315.36 -35.52 315.68 -31.12 ;
      RECT 315.38 -35.545 315.66 -31.12 ;
      RECT 314.7 -21.24 314.98 2.225 ;
      RECT 314.68 -21.24 315 2.2 ;
      RECT 314 -35.52 314.32 2.2 ;
      RECT 314.02 -35.545 314.3 2.2 ;
      RECT 313.34 -35.52 313.62 2.225 ;
      RECT 313.32 -35.52 313.64 2.2 ;
      RECT 312.64 -35.52 312.96 2.2 ;
      RECT 312.66 -35.545 312.94 2.2 ;
      RECT 311.98 -35.52 312.26 2.225 ;
      RECT 311.96 -35.52 312.28 2.2 ;
      RECT 311.28 -35.52 311.6 2.2 ;
      RECT 311.3 -35.545 311.58 2.2 ;
      RECT 310.62 -35.52 310.9 2.225 ;
      RECT 310.6 -35.52 310.92 2.2 ;
      RECT 309.92 -35.52 310.24 2.2 ;
      RECT 309.94 -35.545 310.22 2.2 ;
      RECT 309.26 -24.64 309.54 2.225 ;
      RECT 309.24 -24.64 309.56 2.2 ;
      RECT 308.04 -35.475 308.36 -30.11 ;
      RECT 308.06 -35.495 308.34 -30.11 ;
      RECT 307.9 -20.56 308.18 2.225 ;
      RECT 307.88 -20.56 308.2 2.2 ;
      RECT 306.54 -35.52 306.82 2.225 ;
      RECT 306.52 -35.52 306.84 2.2 ;
      RECT 305.18 -25.32 305.46 2.225 ;
      RECT 305.16 -25.32 305.48 2.2 ;
      RECT 303.82 -17.16 304.1 2.225 ;
      RECT 303.8 -17.16 304.12 2.2 ;
      RECT 302.46 -18.52 302.74 2.225 ;
      RECT 302.44 -18.52 302.76 2.2 ;
      RECT 301.1 -18.52 301.38 2.225 ;
      RECT 301.08 -18.52 301.4 2.2 ;
      RECT 300.4 -35.52 300.72 -31.12 ;
      RECT 300.42 -35.545 300.7 -31.12 ;
      RECT 299.74 -21.24 300.02 2.225 ;
      RECT 299.72 -21.24 300.04 2.2 ;
      RECT 299.04 -35.52 299.36 2.2 ;
      RECT 299.06 -35.545 299.34 2.2 ;
      RECT 298.38 -35.52 298.66 2.225 ;
      RECT 298.36 -35.52 298.68 2.2 ;
      RECT 297.68 -35.52 298 2.2 ;
      RECT 297.7 -35.545 297.98 2.2 ;
      RECT 297.02 -35.52 297.3 2.225 ;
      RECT 297 -35.52 297.32 2.2 ;
      RECT 296.32 -35.52 296.64 2.2 ;
      RECT 296.34 -35.545 296.62 2.2 ;
      RECT 295.66 -35.52 295.94 2.225 ;
      RECT 295.64 -35.52 295.96 2.2 ;
      RECT 294.96 -35.52 295.28 2.2 ;
      RECT 294.98 -35.545 295.26 2.2 ;
      RECT 294.3 -24.64 294.58 2.225 ;
      RECT 294.28 -24.64 294.6 2.2 ;
      RECT 293.14 -35.475 293.46 -30.11 ;
      RECT 293.16 -35.495 293.44 -30.11 ;
      RECT 292.94 -20.56 293.22 2.225 ;
      RECT 292.92 -20.56 293.24 2.2 ;
      RECT 291.58 -35.52 291.86 2.225 ;
      RECT 291.56 -35.52 291.88 2.2 ;
      RECT 290.22 -25.32 290.5 2.225 ;
      RECT 290.2 -25.32 290.52 2.2 ;
      RECT 288.86 -17.16 289.14 2.225 ;
      RECT 288.84 -17.16 289.16 2.2 ;
      RECT 287.5 -18.52 287.78 2.225 ;
      RECT 287.48 -18.52 287.8 2.2 ;
      RECT 286.14 -18.52 286.42 2.225 ;
      RECT 286.12 -18.52 286.44 2.2 ;
      RECT 285.44 -35.52 285.76 -31.12 ;
      RECT 285.46 -35.545 285.74 -31.12 ;
      RECT 284.78 -35.52 285.06 2.225 ;
      RECT 284.76 -35.52 285.08 2.2 ;
      RECT 284.08 -35.52 284.4 2.2 ;
      RECT 284.1 -35.545 284.38 2.2 ;
      RECT 283.42 -35.52 283.7 2.225 ;
      RECT 283.4 -35.52 283.72 2.2 ;
      RECT 282.72 -35.52 283.04 2.2 ;
      RECT 282.74 -35.545 283.02 2.2 ;
      RECT 282.06 -35.52 282.34 2.225 ;
      RECT 282.04 -35.52 282.36 2.2 ;
      RECT 281.36 -35.52 281.68 2.2 ;
      RECT 281.38 -35.545 281.66 2.2 ;
      RECT 280.7 -35.52 280.98 2.225 ;
      RECT 280.68 -35.52 281 2.2 ;
      RECT 280 -35.52 280.32 2.2 ;
      RECT 280.02 -35.545 280.3 2.2 ;
      RECT 279.34 -24.64 279.62 2.225 ;
      RECT 279.32 -24.64 279.64 2.2 ;
      RECT 278.24 -35.475 278.56 -30.11 ;
      RECT 278.26 -35.495 278.54 -30.11 ;
      RECT 277.98 -20.56 278.26 2.225 ;
      RECT 277.96 -20.56 278.28 2.2 ;
      RECT 276.62 -35.52 276.9 2.225 ;
      RECT 276.6 -35.52 276.92 2.2 ;
      RECT 275.26 -25.32 275.54 2.225 ;
      RECT 275.24 -25.32 275.56 2.2 ;
      RECT 273.9 -17.16 274.18 2.225 ;
      RECT 273.88 -17.16 274.2 2.2 ;
      RECT 272.54 -21.92 272.82 2.225 ;
      RECT 272.52 -21.92 272.84 2.2 ;
      RECT 271.18 -18.52 271.46 2.225 ;
      RECT 271.16 -18.52 271.48 2.2 ;
      RECT 270.48 -35.52 270.8 -31.12 ;
      RECT 270.5 -35.545 270.78 -31.12 ;
      RECT 269.82 -35.52 270.1 2.225 ;
      RECT 269.8 -35.52 270.12 2.2 ;
      RECT 269.12 -35.52 269.44 2.2 ;
      RECT 269.14 -35.545 269.42 2.2 ;
      RECT 268.46 -35.52 268.74 2.225 ;
      RECT 268.44 -35.52 268.76 2.2 ;
      RECT 267.76 -35.52 268.08 2.2 ;
      RECT 267.78 -35.545 268.06 2.2 ;
      RECT 267.1 -35.52 267.38 2.225 ;
      RECT 267.08 -35.52 267.4 2.2 ;
      RECT 266.4 -35.52 266.72 2.2 ;
      RECT 266.42 -35.545 266.7 2.2 ;
      RECT 265.74 -35.52 266.02 2.225 ;
      RECT 265.72 -35.52 266.04 2.2 ;
      RECT 265.04 -35.52 265.36 2.2 ;
      RECT 265.06 -35.545 265.34 2.2 ;
      RECT 264.38 -24.64 264.66 2.225 ;
      RECT 264.36 -24.64 264.68 2.2 ;
      RECT 263.34 -35.475 263.66 -30.11 ;
      RECT 263.36 -35.495 263.64 -30.11 ;
      RECT 263.02 -20.56 263.3 2.225 ;
      RECT 263 -20.56 263.32 2.2 ;
      RECT 261.66 -35.52 261.94 2.225 ;
      RECT 261.64 -35.52 261.96 2.2 ;
      RECT 260.3 -25.32 260.58 2.225 ;
      RECT 260.28 -25.32 260.6 2.2 ;
      RECT 258.94 -17.16 259.22 2.225 ;
      RECT 258.92 -17.16 259.24 2.2 ;
      RECT 257.58 -21.92 257.86 2.225 ;
      RECT 257.56 -21.92 257.88 2.2 ;
      RECT 256.22 -18.52 256.5 2.225 ;
      RECT 256.2 -18.52 256.52 2.2 ;
      RECT 255.52 -35.52 255.84 -31.12 ;
      RECT 255.54 -35.545 255.82 -31.12 ;
      RECT 254.86 -35.52 255.14 2.225 ;
      RECT 254.84 -35.52 255.16 2.2 ;
      RECT 254.16 -35.52 254.48 2.2 ;
      RECT 254.18 -35.545 254.46 2.2 ;
      RECT 253.5 -35.52 253.78 2.225 ;
      RECT 253.48 -35.52 253.8 2.2 ;
      RECT 252.8 -35.52 253.12 2.2 ;
      RECT 252.82 -35.545 253.1 2.2 ;
      RECT 252.14 -35.52 252.42 2.225 ;
      RECT 252.12 -35.52 252.44 2.2 ;
      RECT 251.44 -35.52 251.76 2.2 ;
      RECT 251.46 -35.545 251.74 2.2 ;
      RECT 250.78 -35.52 251.06 2.225 ;
      RECT 250.76 -35.52 251.08 2.2 ;
      RECT 250.08 -35.52 250.4 2.2 ;
      RECT 250.1 -35.545 250.38 2.2 ;
      RECT 249.42 -24.64 249.7 2.225 ;
      RECT 249.4 -24.64 249.72 2.2 ;
      RECT 248.44 -35.475 248.76 -30.11 ;
      RECT 248.46 -35.495 248.74 -30.11 ;
      RECT 248.06 -20.56 248.34 2.225 ;
      RECT 248.04 -20.56 248.36 2.2 ;
      RECT 246.7 -35.52 246.98 2.225 ;
      RECT 246.68 -35.52 247 2.2 ;
      RECT 245.34 -17.16 245.62 2.225 ;
      RECT 245.32 -17.16 245.64 2.2 ;
      RECT 243.98 -17.84 244.26 2.225 ;
      RECT 243.96 -17.84 244.28 2.2 ;
      RECT 242.62 -21.92 242.9 2.225 ;
      RECT 242.6 -21.92 242.92 2.2 ;
      RECT 241.26 -18.52 241.54 2.225 ;
      RECT 241.24 -18.52 241.56 2.2 ;
      RECT 240.56 -35.52 240.88 -31.12 ;
      RECT 240.58 -35.545 240.86 -31.12 ;
      RECT 239.9 -35.52 240.18 2.225 ;
      RECT 239.88 -35.52 240.2 2.2 ;
      RECT 239.2 -35.52 239.52 2.2 ;
      RECT 239.22 -35.545 239.5 2.2 ;
      RECT 238.54 -35.52 238.82 2.225 ;
      RECT 238.52 -35.52 238.84 2.2 ;
      RECT 237.84 -35.52 238.16 2.2 ;
      RECT 237.86 -35.545 238.14 2.2 ;
      RECT 237.18 -35.52 237.46 2.225 ;
      RECT 237.16 -35.52 237.48 2.2 ;
      RECT 236.48 -35.52 236.8 2.2 ;
      RECT 236.5 -35.545 236.78 2.2 ;
      RECT 235.82 -35.52 236.1 2.225 ;
      RECT 235.8 -35.52 236.12 2.2 ;
      RECT 235.12 -35.52 235.44 2.2 ;
      RECT 235.14 -35.545 235.42 2.2 ;
      RECT 234.46 -24.64 234.74 2.225 ;
      RECT 234.44 -24.64 234.76 2.2 ;
      RECT 233.54 -35.475 233.86 -30.11 ;
      RECT 233.56 -35.495 233.84 -30.11 ;
      RECT 233.1 -20.56 233.38 2.225 ;
      RECT 233.08 -20.56 233.4 2.2 ;
      RECT 231.74 -35.52 232.02 2.225 ;
      RECT 231.72 -35.52 232.04 2.2 ;
      RECT 230.38 -17.16 230.66 2.225 ;
      RECT 230.36 -17.16 230.68 2.2 ;
      RECT 229.02 -17.84 229.3 2.225 ;
      RECT 229 -17.84 229.32 2.2 ;
      RECT 227.66 -21.92 227.94 2.225 ;
      RECT 227.64 -21.92 227.96 2.2 ;
      RECT 226.3 -18.52 226.58 2.225 ;
      RECT 226.28 -18.52 226.6 2.2 ;
      RECT 225.6 -35.52 225.92 -31.12 ;
      RECT 225.62 -35.545 225.9 -31.12 ;
      RECT 224.94 -35.52 225.22 2.225 ;
      RECT 224.92 -35.52 225.24 2.2 ;
      RECT 224.24 -35.52 224.56 2.2 ;
      RECT 224.26 -35.545 224.54 2.2 ;
      RECT 223.58 -35.52 223.86 2.225 ;
      RECT 223.56 -35.52 223.88 2.2 ;
      RECT 222.88 -35.52 223.2 2.2 ;
      RECT 222.9 -35.545 223.18 2.2 ;
      RECT 222.22 -35.52 222.5 2.225 ;
      RECT 222.2 -35.52 222.52 2.2 ;
      RECT 221.52 -35.52 221.84 2.2 ;
      RECT 221.54 -35.545 221.82 2.2 ;
      RECT 220.86 -35.52 221.14 2.225 ;
      RECT 220.84 -35.52 221.16 2.2 ;
      RECT 220.16 -35.52 220.48 2.2 ;
      RECT 220.18 -35.545 220.46 2.2 ;
      RECT 219.5 -24.64 219.78 2.225 ;
      RECT 219.48 -24.64 219.8 2.2 ;
      RECT 218.64 -35.475 218.96 -30.11 ;
      RECT 218.66 -35.495 218.94 -30.11 ;
      RECT 218.14 -20.56 218.42 2.225 ;
      RECT 218.12 -20.56 218.44 2.2 ;
      RECT 216.78 -25.32 217.06 2.225 ;
      RECT 216.76 -25.32 217.08 2.2 ;
      RECT 215.42 -17.16 215.7 2.225 ;
      RECT 215.4 -17.16 215.72 2.2 ;
      RECT 214.06 -17.84 214.34 2.225 ;
      RECT 214.04 -17.84 214.36 2.2 ;
      RECT 212.7 -21.92 212.98 2.225 ;
      RECT 212.68 -21.92 213 2.2 ;
      RECT 211.34 -18.52 211.62 2.225 ;
      RECT 211.32 -18.52 211.64 2.2 ;
      RECT 210.64 -35.52 210.96 -31.12 ;
      RECT 210.66 -35.545 210.94 -31.12 ;
      RECT 209.98 -35.52 210.26 2.225 ;
      RECT 209.96 -35.52 210.28 2.2 ;
      RECT 209.28 -35.52 209.6 2.2 ;
      RECT 209.3 -35.545 209.58 2.2 ;
      RECT 208.62 -35.52 208.9 2.225 ;
      RECT 208.6 -35.52 208.92 2.2 ;
      RECT 207.92 -35.52 208.24 2.2 ;
      RECT 207.94 -35.545 208.22 2.2 ;
      RECT 207.26 -35.52 207.54 2.225 ;
      RECT 207.24 -35.52 207.56 2.2 ;
      RECT 206.56 -35.52 206.88 2.2 ;
      RECT 206.58 -35.545 206.86 2.2 ;
      RECT 205.9 -35.52 206.18 2.225 ;
      RECT 205.88 -35.52 206.2 2.2 ;
      RECT 205.2 -35.52 205.52 2.2 ;
      RECT 205.22 -35.545 205.5 2.2 ;
      RECT 204.54 -24.64 204.82 2.225 ;
      RECT 204.52 -24.64 204.84 2.2 ;
      RECT 203.74 -35.475 204.06 -30.11 ;
      RECT 203.76 -35.495 204.04 -30.11 ;
      RECT 203.18 -20.56 203.46 2.225 ;
      RECT 203.16 -20.56 203.48 2.2 ;
      RECT 201.82 -25.32 202.1 2.225 ;
      RECT 201.8 -25.32 202.12 2.2 ;
      RECT 200.46 -17.16 200.74 2.225 ;
      RECT 200.44 -17.16 200.76 2.2 ;
      RECT 199.1 -17.84 199.38 2.225 ;
      RECT 199.08 -17.84 199.4 2.2 ;
      RECT 197.74 -21.92 198.02 2.225 ;
      RECT 197.72 -21.92 198.04 2.2 ;
      RECT 196.38 -18.52 196.66 2.225 ;
      RECT 196.36 -18.52 196.68 2.2 ;
      RECT 195.68 -35.52 196 -31.12 ;
      RECT 195.7 -35.545 195.98 -31.12 ;
      RECT 195.02 -35.52 195.3 2.225 ;
      RECT 195 -35.52 195.32 2.2 ;
      RECT 194.32 -35.52 194.64 2.2 ;
      RECT 194.34 -35.545 194.62 2.2 ;
      RECT 193.66 -35.52 193.94 2.225 ;
      RECT 193.64 -35.52 193.96 2.2 ;
      RECT 192.96 -35.52 193.28 2.2 ;
      RECT 192.98 -35.545 193.26 2.2 ;
      RECT 192.3 -35.52 192.58 2.225 ;
      RECT 192.28 -35.52 192.6 2.2 ;
      RECT 191.6 -35.52 191.92 2.2 ;
      RECT 191.62 -35.545 191.9 2.2 ;
      RECT 190.94 -35.52 191.22 2.225 ;
      RECT 190.92 -35.52 191.24 2.2 ;
      RECT 190.24 -35.52 190.56 2.2 ;
      RECT 190.26 -35.545 190.54 2.2 ;
      RECT 189.58 -24.64 189.86 2.225 ;
      RECT 189.56 -24.64 189.88 2.2 ;
      RECT 188.84 -35.475 189.16 -30.11 ;
      RECT 188.86 -35.495 189.14 -30.11 ;
      RECT 188.22 -20.56 188.5 2.225 ;
      RECT 188.2 -20.56 188.52 2.2 ;
      RECT 186.86 -25.32 187.14 2.225 ;
      RECT 186.84 -25.32 187.16 2.2 ;
      RECT 185.5 -17.16 185.78 2.225 ;
      RECT 185.48 -17.16 185.8 2.2 ;
      RECT 184.14 -17.84 184.42 2.225 ;
      RECT 184.12 -17.84 184.44 2.2 ;
      RECT 182.78 -21.92 183.06 2.225 ;
      RECT 182.76 -21.92 183.08 2.2 ;
      RECT 181.42 -18.52 181.7 2.225 ;
      RECT 181.4 -18.52 181.72 2.2 ;
      RECT 180.72 -35.52 181.04 -31.12 ;
      RECT 180.74 -35.545 181.02 -31.12 ;
      RECT 180.06 -35.52 180.34 2.225 ;
      RECT 180.04 -35.52 180.36 2.2 ;
      RECT 179.36 -35.52 179.68 2.2 ;
      RECT 179.38 -35.545 179.66 2.2 ;
      RECT 178.7 -35.52 178.98 2.225 ;
      RECT 178.68 -35.52 179 2.2 ;
      RECT 178 -35.52 178.32 2.2 ;
      RECT 178.02 -35.545 178.3 2.2 ;
      RECT 177.34 -35.52 177.62 2.225 ;
      RECT 177.32 -35.52 177.64 2.2 ;
      RECT 176.64 -35.52 176.96 2.2 ;
      RECT 176.66 -35.545 176.94 2.2 ;
      RECT 175.98 -35.52 176.26 2.225 ;
      RECT 175.96 -35.52 176.28 2.2 ;
      RECT 175.28 -35.52 175.6 2.2 ;
      RECT 175.3 -35.545 175.58 2.2 ;
      RECT 174.62 -20.56 174.9 2.225 ;
      RECT 174.6 -20.56 174.92 2.2 ;
      RECT 173.94 -35.475 174.26 -30.11 ;
      RECT 173.96 -35.495 174.24 -30.11 ;
      RECT 173.26 -21.24 173.54 2.225 ;
      RECT 173.24 -21.24 173.56 2.2 ;
      RECT 171.9 -25.32 172.18 2.225 ;
      RECT 171.88 -25.32 172.2 2.2 ;
      RECT 170.54 -17.16 170.82 2.225 ;
      RECT 170.52 -17.16 170.84 2.2 ;
      RECT 169.18 -17.84 169.46 2.225 ;
      RECT 169.16 -17.84 169.48 2.2 ;
      RECT 167.82 -21.92 168.1 2.225 ;
      RECT 167.8 -21.92 168.12 2.2 ;
      RECT 166.46 -18.52 166.74 2.225 ;
      RECT 166.44 -18.52 166.76 2.2 ;
      RECT 165.76 -35.52 166.08 -31.12 ;
      RECT 165.78 -35.545 166.06 -31.12 ;
      RECT 165.1 -35.52 165.38 2.225 ;
      RECT 165.08 -35.52 165.4 2.2 ;
      RECT 164.4 -35.52 164.72 2.2 ;
      RECT 164.42 -35.545 164.7 2.2 ;
      RECT 163.74 -35.52 164.02 2.225 ;
      RECT 163.72 -35.52 164.04 2.2 ;
      RECT 163.04 -35.52 163.36 2.2 ;
      RECT 163.06 -35.545 163.34 2.2 ;
      RECT 162.38 -35.52 162.66 2.225 ;
      RECT 162.36 -35.52 162.68 2.2 ;
      RECT 161.68 -35.52 162 2.2 ;
      RECT 161.7 -35.545 161.98 2.2 ;
      RECT 161.02 -35.52 161.3 2.225 ;
      RECT 161 -35.52 161.32 2.2 ;
      RECT 159.66 -20.56 159.94 2.225 ;
      RECT 159.64 -20.56 159.96 2.2 ;
      RECT 159.04 -35.475 159.36 -30.11 ;
      RECT 159.06 -35.495 159.34 -30.11 ;
      RECT 158.3 -21.24 158.58 2.225 ;
      RECT 158.28 -21.24 158.6 2.2 ;
      RECT 156.94 -25.32 157.22 2.225 ;
      RECT 156.92 -25.32 157.24 2.2 ;
      RECT 155.58 -17.16 155.86 2.225 ;
      RECT 155.56 -17.16 155.88 2.2 ;
      RECT 154.22 -17.84 154.5 2.225 ;
      RECT 154.2 -17.84 154.52 2.2 ;
      RECT 152.86 -21.92 153.14 2.225 ;
      RECT 152.84 -21.92 153.16 2.2 ;
      RECT 151.5 -18.52 151.78 2.225 ;
      RECT 151.48 -18.52 151.8 2.2 ;
      RECT 150.8 -35.52 151.12 -31.12 ;
      RECT 150.82 -35.545 151.1 -31.12 ;
      RECT 150.14 -35.52 150.42 2.225 ;
      RECT 150.12 -35.52 150.44 2.2 ;
      RECT 149.44 -35.52 149.76 2.2 ;
      RECT 149.46 -35.545 149.74 2.2 ;
      RECT 148.78 -35.52 149.06 2.225 ;
      RECT 148.76 -35.52 149.08 2.2 ;
      RECT 148.08 -35.52 148.4 2.2 ;
      RECT 148.1 -35.545 148.38 2.2 ;
      RECT 147.42 -35.52 147.7 2.225 ;
      RECT 147.4 -35.52 147.72 2.2 ;
      RECT 146.72 -35.52 147.04 2.2 ;
      RECT 146.74 -35.545 147.02 2.2 ;
      RECT 146.06 -35.52 146.34 2.225 ;
      RECT 146.04 -35.52 146.36 2.2 ;
      RECT 144.7 -20.56 144.98 2.225 ;
      RECT 144.68 -20.56 145 2.2 ;
      RECT 144.14 -35.475 144.46 -30.11 ;
      RECT 144.16 -35.495 144.44 -30.11 ;
      RECT 143.34 -21.24 143.62 2.225 ;
      RECT 143.32 -21.24 143.64 2.2 ;
      RECT 141.98 -25.32 142.26 2.225 ;
      RECT 141.96 -25.32 142.28 2.2 ;
      RECT 140.62 -17.16 140.9 2.225 ;
      RECT 140.6 -17.16 140.92 2.2 ;
      RECT 139.26 -17.84 139.54 2.225 ;
      RECT 139.24 -17.84 139.56 2.2 ;
      RECT 137.9 -18.52 138.18 2.225 ;
      RECT 137.88 -18.52 138.2 2.2 ;
      RECT 136.54 -21.24 136.82 2.225 ;
      RECT 136.52 -21.24 136.84 2.2 ;
      RECT 135.84 -35.52 136.16 -31.12 ;
      RECT 135.86 -35.545 136.14 -31.12 ;
      RECT 135.18 -35.52 135.46 2.225 ;
      RECT 135.16 -35.52 135.48 2.2 ;
      RECT 134.48 -35.52 134.8 2.2 ;
      RECT 134.5 -35.545 134.78 2.2 ;
      RECT 133.82 -35.52 134.1 2.225 ;
      RECT 133.8 -35.52 134.12 2.2 ;
      RECT 133.12 -35.52 133.44 2.2 ;
      RECT 133.14 -35.545 133.42 2.2 ;
      RECT 132.46 -35.52 132.74 2.225 ;
      RECT 132.44 -35.52 132.76 2.2 ;
      RECT 131.76 -35.52 132.08 2.2 ;
      RECT 131.78 -35.545 132.06 2.2 ;
      RECT 131.1 -35.52 131.38 2.225 ;
      RECT 131.08 -35.52 131.4 2.2 ;
      RECT 129.74 -20.56 130.02 2.225 ;
      RECT 129.72 -20.56 130.04 2.2 ;
      RECT 129.24 -35.475 129.56 -30.11 ;
      RECT 129.26 -35.495 129.54 -30.11 ;
      RECT 128.38 -21.24 128.66 2.225 ;
      RECT 128.36 -21.24 128.68 2.2 ;
      RECT 127.02 -25.32 127.3 2.225 ;
      RECT 127 -25.32 127.32 2.2 ;
      RECT 125.66 -17.16 125.94 2.225 ;
      RECT 125.64 -17.16 125.96 2.2 ;
      RECT 124.3 -17.84 124.58 2.225 ;
      RECT 124.28 -17.84 124.6 2.2 ;
      RECT 122.94 -18.52 123.22 2.225 ;
      RECT 122.92 -18.52 123.24 2.2 ;
      RECT 122.24 -35.52 122.56 -31.12 ;
      RECT 122.26 -35.545 122.54 -31.12 ;
      RECT 121.58 -21.24 121.86 2.225 ;
      RECT 121.56 -21.24 121.88 2.2 ;
      RECT 120.88 -35.52 121.2 2.2 ;
      RECT 120.9 -35.545 121.18 2.2 ;
      RECT 120.22 -35.52 120.5 2.225 ;
      RECT 120.2 -35.52 120.52 2.2 ;
      RECT 119.52 -35.52 119.84 2.2 ;
      RECT 119.54 -35.545 119.82 2.2 ;
      RECT 118.86 -35.52 119.14 2.225 ;
      RECT 118.84 -35.52 119.16 2.2 ;
      RECT 118.16 -35.52 118.48 2.2 ;
      RECT 118.18 -35.545 118.46 2.2 ;
      RECT 117.5 -35.52 117.78 2.225 ;
      RECT 117.48 -35.52 117.8 2.2 ;
      RECT 116.8 -35.52 117.12 2.2 ;
      RECT 116.82 -35.545 117.1 2.2 ;
      RECT 116.14 -35.52 116.42 2.225 ;
      RECT 116.12 -35.52 116.44 2.2 ;
      RECT 114.78 -20.56 115.06 2.225 ;
      RECT 114.76 -20.56 115.08 2.2 ;
      RECT 114.34 -35.475 114.66 -30.11 ;
      RECT 114.36 -35.495 114.64 -30.11 ;
      RECT 113.42 -21.24 113.7 2.225 ;
      RECT 113.4 -21.24 113.72 2.2 ;
      RECT 112.06 -25.32 112.34 2.225 ;
      RECT 112.04 -25.32 112.36 2.2 ;
      RECT 110.7 -17.16 110.98 2.225 ;
      RECT 110.68 -17.16 111 2.2 ;
      RECT 109.34 -17.84 109.62 2.225 ;
      RECT 109.32 -17.84 109.64 2.2 ;
      RECT 107.98 -18.52 108.26 2.225 ;
      RECT 107.96 -18.52 108.28 2.2 ;
      RECT 107.28 -35.52 107.6 -31.12 ;
      RECT 107.3 -35.545 107.58 -31.12 ;
      RECT 106.62 -21.24 106.9 2.225 ;
      RECT 106.6 -21.24 106.92 2.2 ;
      RECT 105.92 -35.52 106.24 2.2 ;
      RECT 105.94 -35.545 106.22 2.2 ;
      RECT 105.26 -35.52 105.54 2.225 ;
      RECT 105.24 -35.52 105.56 2.2 ;
      RECT 104.56 -35.52 104.88 2.2 ;
      RECT 104.58 -35.545 104.86 2.2 ;
      RECT 103.9 -35.52 104.18 2.225 ;
      RECT 103.88 -35.52 104.2 2.2 ;
      RECT 103.2 -35.52 103.52 2.2 ;
      RECT 103.22 -35.545 103.5 2.2 ;
      RECT 102.54 -35.52 102.82 2.225 ;
      RECT 102.52 -35.52 102.84 2.2 ;
      RECT 101.84 -35.52 102.16 2.2 ;
      RECT 101.86 -35.545 102.14 2.2 ;
      RECT 101.18 -35.52 101.46 2.225 ;
      RECT 101.16 -35.52 101.48 2.2 ;
      RECT 99.82 -20.56 100.1 2.225 ;
      RECT 99.8 -20.56 100.12 2.2 ;
      RECT 99.44 -35.475 99.76 -30.11 ;
      RECT 99.46 -35.495 99.74 -30.11 ;
      RECT 98.46 -21.24 98.74 2.225 ;
      RECT 98.44 -21.24 98.76 2.2 ;
      RECT 97.1 -25.32 97.38 2.225 ;
      RECT 97.08 -25.32 97.4 2.2 ;
      RECT 95.74 -17.16 96.02 2.225 ;
      RECT 95.72 -17.16 96.04 2.2 ;
      RECT 94.38 -17.84 94.66 2.225 ;
      RECT 94.36 -17.84 94.68 2.2 ;
      RECT 93.02 -18.52 93.3 2.225 ;
      RECT 93 -18.52 93.32 2.2 ;
      RECT 92.32 -35.52 92.64 -31.12 ;
      RECT 92.34 -35.545 92.62 -31.12 ;
      RECT 91.66 -21.24 91.94 2.225 ;
      RECT 91.64 -21.24 91.96 2.2 ;
      RECT 90.96 -35.52 91.28 2.2 ;
      RECT 90.98 -35.545 91.26 2.2 ;
      RECT 90.3 -35.52 90.58 2.225 ;
      RECT 90.28 -35.52 90.6 2.2 ;
      RECT 89.6 -35.52 89.92 2.2 ;
      RECT 89.62 -35.545 89.9 2.2 ;
      RECT 88.94 -35.52 89.22 2.225 ;
      RECT 88.92 -35.52 89.24 2.2 ;
      RECT 88.24 -35.52 88.56 2.2 ;
      RECT 88.26 -35.545 88.54 2.2 ;
      RECT 87.58 -35.52 87.86 2.225 ;
      RECT 87.56 -35.52 87.88 2.2 ;
      RECT 86.88 -35.52 87.2 2.2 ;
      RECT 86.9 -35.545 87.18 2.2 ;
      RECT 86.22 -35.52 86.5 2.225 ;
      RECT 86.2 -35.52 86.52 2.2 ;
      RECT 84.86 -20.56 85.14 2.225 ;
      RECT 84.84 -20.56 85.16 2.2 ;
      RECT 84.54 -35.475 84.86 -30.11 ;
      RECT 84.56 -35.495 84.84 -30.11 ;
      RECT 83.5 -21.24 83.78 2.225 ;
      RECT 83.48 -21.24 83.8 2.2 ;
      RECT 82.14 -25.32 82.42 2.225 ;
      RECT 82.12 -25.32 82.44 2.2 ;
      RECT 80.78 -17.16 81.06 2.225 ;
      RECT 80.76 -17.16 81.08 2.2 ;
      RECT 79.42 -18.52 79.7 2.225 ;
      RECT 79.4 -18.52 79.72 2.2 ;
      RECT 78.06 -18.52 78.34 2.225 ;
      RECT 78.04 -18.52 78.36 2.2 ;
      RECT 77.36 -35.52 77.68 -31.12 ;
      RECT 77.38 -35.545 77.66 -31.12 ;
      RECT 76.7 -21.24 76.98 2.225 ;
      RECT 76.68 -21.24 77 2.2 ;
      RECT 76 -35.52 76.32 2.2 ;
      RECT 76.02 -35.545 76.3 2.2 ;
      RECT 75.34 -35.52 75.62 2.225 ;
      RECT 75.32 -35.52 75.64 2.2 ;
      RECT 74.64 -35.52 74.96 2.2 ;
      RECT 74.66 -35.545 74.94 2.2 ;
      RECT 73.98 -35.52 74.26 2.225 ;
      RECT 73.96 -35.52 74.28 2.2 ;
      RECT 73.28 -35.52 73.6 2.2 ;
      RECT 73.3 -35.545 73.58 2.2 ;
      RECT 72.62 -35.52 72.9 2.225 ;
      RECT 72.6 -35.52 72.92 2.2 ;
      RECT 71.92 -35.52 72.24 2.2 ;
      RECT 71.94 -35.545 72.22 2.2 ;
      RECT 71.26 -35.52 71.54 2.225 ;
      RECT 71.24 -35.52 71.56 2.2 ;
      RECT 69.9 -20.56 70.18 2.225 ;
      RECT 69.88 -20.56 70.2 2.2 ;
      RECT 69.64 -35.475 69.96 -30.11 ;
      RECT 69.66 -35.495 69.94 -30.11 ;
      RECT 68.54 -21.24 68.82 2.225 ;
      RECT 68.52 -21.24 68.84 2.2 ;
      RECT 67.18 -25.32 67.46 2.225 ;
      RECT 67.16 -25.32 67.48 2.2 ;
      RECT 65.82 -17.16 66.1 2.225 ;
      RECT 65.8 -17.16 66.12 2.2 ;
      RECT 64.46 -18.52 64.74 2.225 ;
      RECT 64.44 -18.52 64.76 2.2 ;
      RECT 63.1 -18.52 63.38 2.225 ;
      RECT 63.08 -18.52 63.4 2.2 ;
      RECT 62.4 -35.52 62.72 -31.12 ;
      RECT 62.42 -35.545 62.7 -31.12 ;
      RECT 61.74 -21.24 62.02 2.225 ;
      RECT 61.72 -21.24 62.04 2.2 ;
      RECT 61.04 -35.52 61.36 2.2 ;
      RECT 61.06 -35.545 61.34 2.2 ;
      RECT 60.38 -35.52 60.66 2.225 ;
      RECT 60.36 -35.52 60.68 2.2 ;
      RECT 59.68 -35.52 60 2.2 ;
      RECT 59.7 -35.545 59.98 2.2 ;
      RECT 59.02 -35.52 59.3 2.225 ;
      RECT 59 -35.52 59.32 2.2 ;
      RECT 58.32 -35.52 58.64 2.2 ;
      RECT 58.34 -35.545 58.62 2.2 ;
      RECT 57.66 -35.52 57.94 2.225 ;
      RECT 57.64 -35.52 57.96 2.2 ;
      RECT 56.96 -35.52 57.28 2.2 ;
      RECT 56.98 -35.545 57.26 2.2 ;
      RECT 56.3 -35.52 56.58 2.225 ;
      RECT 56.28 -35.52 56.6 2.2 ;
      RECT 54.94 -20.56 55.22 2.225 ;
      RECT 54.92 -20.56 55.24 2.2 ;
      RECT 54.74 -35.475 55.06 -30.11 ;
      RECT 54.76 -35.495 55.04 -30.11 ;
      RECT 53.58 -21.24 53.86 2.225 ;
      RECT 53.56 -21.24 53.88 2.2 ;
      RECT 52.22 -25.32 52.5 2.225 ;
      RECT 52.2 -25.32 52.52 2.2 ;
      RECT 50.86 -17.16 51.14 2.225 ;
      RECT 50.84 -17.16 51.16 2.2 ;
      RECT 49.5 -18.52 49.78 2.225 ;
      RECT 49.48 -18.52 49.8 2.2 ;
      RECT 48.14 -18.52 48.42 2.225 ;
      RECT 48.12 -18.52 48.44 2.2 ;
      RECT 47.44 -35.52 47.76 -31.12 ;
      RECT 47.46 -35.545 47.74 -31.12 ;
      RECT 46.78 -21.24 47.06 2.225 ;
      RECT 46.76 -21.24 47.08 2.2 ;
      RECT 46.08 -35.52 46.4 2.2 ;
      RECT 46.1 -35.545 46.38 2.2 ;
      RECT 45.42 -35.52 45.7 2.225 ;
      RECT 45.4 -35.52 45.72 2.2 ;
      RECT 44.72 -35.52 45.04 2.2 ;
      RECT 44.74 -35.545 45.02 2.2 ;
      RECT 44.06 -35.52 44.34 2.225 ;
      RECT 44.04 -35.52 44.36 2.2 ;
      RECT 43.36 -35.52 43.68 2.2 ;
      RECT 43.38 -35.545 43.66 2.2 ;
      RECT 42.7 -35.52 42.98 2.225 ;
      RECT 42.68 -35.52 43 2.2 ;
      RECT 42 -35.52 42.32 2.2 ;
      RECT 42.02 -35.545 42.3 2.2 ;
      RECT 41.34 -35.52 41.62 2.225 ;
      RECT 41.32 -35.52 41.64 2.2 ;
      RECT 39.98 -20.56 40.26 2.225 ;
      RECT 39.96 -20.56 40.28 2.2 ;
      RECT 39.84 -35.475 40.16 -30.11 ;
      RECT 39.86 -35.495 40.14 -30.11 ;
      RECT 38.62 -21.24 38.9 2.225 ;
      RECT 38.6 -21.24 38.92 2.2 ;
      RECT 37.26 -25.32 37.54 2.225 ;
      RECT 37.24 -25.32 37.56 2.2 ;
      RECT 35.9 -17.16 36.18 2.225 ;
      RECT 35.88 -17.16 36.2 2.2 ;
      RECT 34.54 -18.52 34.82 2.225 ;
      RECT 34.52 -18.52 34.84 2.2 ;
      RECT 33.18 -18.52 33.46 2.225 ;
      RECT 33.16 -18.52 33.48 2.2 ;
      RECT 32.48 -35.52 32.8 -31.12 ;
      RECT 32.5 -35.545 32.78 -31.12 ;
      RECT 31.82 -21.24 32.1 2.225 ;
      RECT 31.8 -21.24 32.12 2.2 ;
      RECT 31.12 -35.52 31.44 2.2 ;
      RECT 31.14 -35.545 31.42 2.2 ;
      RECT 30.46 -35.52 30.74 2.225 ;
      RECT 30.44 -35.52 30.76 2.2 ;
      RECT 29.76 -35.52 30.08 2.2 ;
      RECT 29.78 -35.545 30.06 2.2 ;
      RECT 29.1 -35.52 29.38 2.225 ;
      RECT 29.08 -35.52 29.4 2.2 ;
      RECT 28.4 -35.52 28.72 2.2 ;
      RECT 28.42 -35.545 28.7 2.2 ;
      RECT 27.74 -35.52 28.02 2.225 ;
      RECT 27.72 -35.52 28.04 2.2 ;
      RECT 27.04 -35.52 27.36 2.2 ;
      RECT 27.06 -35.545 27.34 2.2 ;
      RECT 26.38 -35.52 26.66 2.225 ;
      RECT 26.36 -35.52 26.68 2.2 ;
      RECT 25.02 -20.56 25.3 2.225 ;
      RECT 25 -20.56 25.32 2.2 ;
      RECT 24.94 -35.475 25.26 -30.11 ;
      RECT 24.96 -35.495 25.24 -30.11 ;
      RECT 23.66 -21.24 23.94 2.225 ;
      RECT 23.64 -21.24 23.96 2.2 ;
      RECT 22.3 -25.32 22.58 2.225 ;
      RECT 22.28 -25.32 22.6 2.2 ;
      RECT 20.94 -17.16 21.22 2.225 ;
      RECT 20.92 -17.16 21.24 2.2 ;
      RECT 19.58 -18.52 19.86 2.225 ;
      RECT 19.56 -18.52 19.88 2.2 ;
      RECT 18.22 -18.52 18.5 2.225 ;
      RECT 18.2 -18.52 18.52 2.2 ;
      RECT 17.52 -35.52 17.84 -31.12 ;
      RECT 17.54 -35.545 17.82 -31.12 ;
      RECT 16.86 -21.24 17.14 2.225 ;
      RECT 16.84 -21.24 17.16 2.2 ;
      RECT 16.16 -35.52 16.48 2.2 ;
      RECT 16.18 -35.545 16.46 2.2 ;
      RECT 15.5 -35.52 15.78 2.225 ;
      RECT 15.48 -35.52 15.8 2.2 ;
      RECT 14.8 -35.52 15.12 2.2 ;
      RECT 14.82 -35.545 15.1 2.2 ;
      RECT 14.14 -35.52 14.42 2.225 ;
      RECT 14.12 -35.52 14.44 2.2 ;
      RECT 13.44 -35.52 13.76 2.2 ;
      RECT 13.46 -35.545 13.74 2.2 ;
      RECT 12.78 -35.52 13.06 2.225 ;
      RECT 12.76 -35.52 13.08 2.2 ;
      RECT 12.08 -35.52 12.4 2.2 ;
      RECT 12.1 -35.545 12.38 2.2 ;
      RECT 11.42 -35.52 11.7 2.225 ;
      RECT 11.4 -35.52 11.72 2.2 ;
      RECT 10.72 -35.52 11.04 2.2 ;
      RECT 10.74 -35.545 11.02 2.2 ;
      RECT 10.06 -20.56 10.34 2.225 ;
      RECT 10.04 -20.56 10.36 2.2 ;
      RECT 9.41 -35.475 9.73 -25.07 ;
      RECT 9.43 -35.495 9.71 -25.07 ;
      RECT 8.7 -35.52 8.98 2.225 ;
      RECT 8.68 -35.52 9 2.2 ;
      RECT 7.34 -34.16 7.62 2.225 ;
      RECT 7.32 -34.16 7.64 2.2 ;
      RECT 5.98 -17.84 6.26 2.225 ;
      RECT 5.96 -17.84 6.28 2.2 ;
      RECT 5.28 -35.52 5.6 -24.32 ;
      RECT 5.3 -35.545 5.58 -24.32 ;
      RECT 4.62 -18.52 4.9 2.225 ;
      RECT 4.6 -18.52 4.92 2.2 ;
      RECT 3.92 -35.52 4.24 -25 ;
      RECT 3.94 -35.545 4.22 -25 ;
      RECT 3.26 -21.92 3.54 2.225 ;
      RECT 3.24 -21.92 3.56 2.2 ;
      RECT 2.56 -35.52 2.88 -25.68 ;
      RECT 2.58 -35.545 2.86 -25.68 ;
      RECT 1.9 -21.24 2.18 2.225 ;
      RECT 1.88 -21.24 2.2 2.2 ;
      RECT 1.2 -35.52 1.52 2.2 ;
      RECT 1.22 -35.545 1.5 2.2 ;
      RECT 0.54 -35.52 0.82 2.225 ;
      RECT 0.52 -35.52 0.84 2.2 ;
      RECT -0.16 -35.52 0.16 2.2 ;
      RECT -0.14 -35.545 0.14 2.2 ;
      RECT -0.82 -35.52 -0.54 2.225 ;
      RECT -0.84 -35.52 -0.52 2.2 ;
      RECT -1.52 -35.52 -1.2 2.2 ;
      RECT -1.5 -35.545 -1.22 2.2 ;
      RECT 949.12 -20.56 949.44 2.2 ;
      RECT 948.74 -35.47 949.06 -21.29 ;
      RECT 947.76 -21.24 948.08 2.2 ;
      RECT 946.4 -34.16 946.72 2.2 ;
      RECT 945.04 -34.16 945.36 2.2 ;
      RECT 943.68 -18.52 944 2.2 ;
      RECT 943 -35.52 943.32 -25 ;
      RECT 942.32 -18.52 942.64 2.2 ;
      RECT 941.64 -35.52 941.96 -25.68 ;
      RECT 940.96 -21.24 941.28 2.2 ;
      RECT 934.47 -35.47 934.79 -25.07 ;
      RECT 934.16 -20.56 934.48 2.2 ;
      RECT 932.8 -35.52 933.12 -31.12 ;
      RECT 932.8 -21.24 933.12 2.2 ;
      RECT 931.44 -25.32 931.76 2.2 ;
      RECT 931.32 -34.87 931.64 -26.325 ;
      RECT 930.08 -17.16 930.4 2.2 ;
      RECT 928.8 -34.87 929.12 -29.475 ;
      RECT 928.72 -18.52 929.04 2.2 ;
      RECT 927.36 -18.52 927.68 2.2 ;
      RECT 926.68 -35.52 927 -31.12 ;
      RECT 926 -21.24 926.32 2.2 ;
      RECT 919.57 -35.47 919.89 -25.07 ;
      RECT 919.2 -20.56 919.52 2.2 ;
      RECT 917.84 -35.52 918.16 -31.12 ;
      RECT 917.84 -21.24 918.16 2.2 ;
      RECT 916.48 -25.32 916.8 2.2 ;
      RECT 916.42 -34.87 916.74 -26.325 ;
      RECT 915.12 -17.16 915.44 2.2 ;
      RECT 913.9 -34.87 914.22 -29.475 ;
      RECT 913.76 -18.52 914.08 2.2 ;
      RECT 912.4 -18.52 912.72 2.2 ;
      RECT 911.72 -35.52 912.04 -31.12 ;
      RECT 911.04 -21.24 911.36 2.2 ;
      RECT 904.67 -35.47 904.99 -25.07 ;
      RECT 904.24 -20.56 904.56 2.2 ;
      RECT 902.88 -35.52 903.2 -31.12 ;
      RECT 902.88 -21.24 903.2 2.2 ;
      RECT 901.52 -34.87 901.84 -26.325 ;
      RECT 901.52 -25.32 901.84 2.2 ;
      RECT 900.16 -17.16 900.48 2.2 ;
      RECT 899 -34.87 899.32 -29.475 ;
      RECT 898.8 -18.52 899.12 2.2 ;
      RECT 897.44 -18.52 897.76 2.2 ;
      RECT 896.76 -35.52 897.08 -31.12 ;
      RECT 896.08 -21.24 896.4 2.2 ;
      RECT 889.77 -35.47 890.09 -25.07 ;
      RECT 889.28 -20.56 889.6 2.2 ;
      RECT 887.92 -35.52 888.24 -31.12 ;
      RECT 887.92 -21.24 888.24 2.2 ;
      RECT 886.62 -34.87 886.94 -26.325 ;
      RECT 886.56 -25.32 886.88 2.2 ;
      RECT 885.2 -17.16 885.52 2.2 ;
      RECT 884.1 -34.87 884.42 -29.475 ;
      RECT 883.84 -18.52 884.16 2.2 ;
      RECT 882.48 -18.52 882.8 2.2 ;
      RECT 881.8 -35.52 882.12 -31.12 ;
      RECT 881.12 -21.24 881.44 2.2 ;
      RECT 874.87 -35.47 875.19 -25.07 ;
      RECT 874.32 -20.56 874.64 2.2 ;
      RECT 872.96 -35.52 873.28 -31.12 ;
      RECT 872.96 -21.24 873.28 2.2 ;
      RECT 871.72 -34.87 872.04 -26.325 ;
      RECT 871.6 -25.32 871.92 2.2 ;
      RECT 870.24 -17.16 870.56 2.2 ;
      RECT 869.2 -34.87 869.52 -29.475 ;
      RECT 868.88 -18.52 869.2 2.2 ;
      RECT 867.52 -18.52 867.84 2.2 ;
      RECT 866.84 -35.52 867.16 -31.12 ;
      RECT 866.16 -21.24 866.48 2.2 ;
      RECT 859.97 -35.47 860.29 -25.07 ;
      RECT 859.36 -20.56 859.68 2.2 ;
      RECT 858 -35.52 858.32 2.2 ;
      RECT 856.82 -34.87 857.14 -26.325 ;
      RECT 856.64 -25.32 856.96 2.2 ;
      RECT 855.28 -17.16 855.6 2.2 ;
      RECT 854.3 -34.87 854.62 -29.475 ;
      RECT 853.92 -18.52 854.24 2.2 ;
      RECT 852.56 -18.52 852.88 2.2 ;
      RECT 851.88 -35.52 852.2 -31.12 ;
      RECT 851.2 -21.24 851.52 2.2 ;
      RECT 845.07 -35.47 845.39 -25.07 ;
      RECT 844.4 -20.56 844.72 2.2 ;
      RECT 843.72 -35.52 844.04 -31.12 ;
      RECT 843.04 -35.52 843.36 2.2 ;
      RECT 841.92 -34.87 842.24 -26.325 ;
      RECT 841.68 -25.32 842 2.2 ;
      RECT 840.32 -17.16 840.64 2.2 ;
      RECT 839.4 -34.87 839.72 -29.475 ;
      RECT 838.96 -18.52 839.28 2.2 ;
      RECT 837.6 -18.52 837.92 2.2 ;
      RECT 836.92 -35.52 837.24 -31.12 ;
      RECT 836.24 -21.24 836.56 2.2 ;
      RECT 830.8 -24.64 831.12 2.2 ;
      RECT 830.17 -35.47 830.49 -25.07 ;
      RECT 829.44 -20.56 829.76 2.2 ;
      RECT 828.76 -35.52 829.08 -31.12 ;
      RECT 828.08 -35.52 828.4 2.2 ;
      RECT 827.02 -34.87 827.34 -26.325 ;
      RECT 826.72 -25.32 827.04 2.2 ;
      RECT 825.36 -17.16 825.68 2.2 ;
      RECT 824.5 -34.87 824.82 -29.475 ;
      RECT 824 -18.52 824.32 2.2 ;
      RECT 822.64 -18.52 822.96 2.2 ;
      RECT 821.96 -35.52 822.28 -31.12 ;
      RECT 821.28 -21.24 821.6 2.2 ;
      RECT 815.84 -24.64 816.16 2.2 ;
      RECT 815.27 -35.47 815.59 -25.07 ;
      RECT 814.48 -20.56 814.8 2.2 ;
      RECT 813.8 -35.52 814.12 -31.12 ;
      RECT 813.12 -35.52 813.44 2.2 ;
      RECT 812.12 -34.87 812.44 -26.325 ;
      RECT 811.76 -25.32 812.08 2.2 ;
      RECT 810.4 -17.16 810.72 2.2 ;
      RECT 809.6 -34.87 809.92 -29.475 ;
      RECT 809.04 -18.52 809.36 2.2 ;
      RECT 807.68 -18.52 808 2.2 ;
      RECT 807 -35.52 807.32 -31.12 ;
      RECT 806.32 -21.24 806.64 2.2 ;
      RECT 800.88 -24.64 801.2 2.2 ;
      RECT 800.37 -35.47 800.69 -25.07 ;
      RECT 799.52 -20.56 799.84 2.2 ;
      RECT 798.84 -35.52 799.16 -31.12 ;
      RECT 798.16 -35.52 798.48 2.2 ;
      RECT 797.22 -34.87 797.54 -26.325 ;
      RECT 796.8 -25.32 797.12 2.2 ;
      RECT 795.44 -17.16 795.76 2.2 ;
      RECT 794.7 -34.87 795.02 -29.475 ;
      RECT 794.08 -18.52 794.4 2.2 ;
      RECT 792.72 -18.52 793.04 2.2 ;
      RECT 792.04 -35.52 792.36 -31.12 ;
      RECT 785.92 -24.64 786.24 2.2 ;
      RECT 785.47 -35.47 785.79 -25.07 ;
      RECT 784.56 -20.56 784.88 2.2 ;
      RECT 783.88 -35.52 784.2 -31.12 ;
      RECT 783.2 -35.52 783.52 2.2 ;
      RECT 782.32 -34.87 782.64 -26.325 ;
      RECT 781.84 -25.32 782.16 2.2 ;
      RECT 780.48 -17.16 780.8 2.2 ;
      RECT 779.8 -34.87 780.12 -29.475 ;
      RECT 779.12 -21.92 779.44 2.2 ;
      RECT 777.76 -18.52 778.08 2.2 ;
      RECT 777.08 -35.52 777.4 -31.12 ;
      RECT 770.96 -24.64 771.28 2.2 ;
      RECT 770.57 -35.47 770.89 -25.07 ;
      RECT 769.6 -20.56 769.92 2.2 ;
      RECT 768.92 -35.52 769.24 -31.12 ;
      RECT 768.24 -35.52 768.56 2.2 ;
      RECT 767.42 -34.87 767.74 -26.325 ;
      RECT 766.88 -25.32 767.2 2.2 ;
      RECT 765.52 -17.16 765.84 2.2 ;
      RECT 764.9 -34.87 765.22 -29.475 ;
      RECT 764.16 -21.92 764.48 2.2 ;
      RECT 762.8 -18.52 763.12 2.2 ;
      RECT 762.12 -35.52 762.44 -31.12 ;
      RECT 756 -24.64 756.32 2.2 ;
      RECT 755.67 -35.47 755.99 -25.07 ;
      RECT 754.64 -20.56 754.96 2.2 ;
      RECT 753.96 -35.52 754.28 -31.12 ;
      RECT 753.28 -35.52 753.6 2.2 ;
      RECT 752.52 -34.87 752.84 -26.325 ;
      RECT 751.92 -17.16 752.24 2.2 ;
      RECT 750.56 -17.84 750.88 2.2 ;
      RECT 750 -34.87 750.32 -29.475 ;
      RECT 749.2 -21.92 749.52 2.2 ;
      RECT 747.84 -18.52 748.16 2.2 ;
      RECT 747.16 -35.52 747.48 -31.12 ;
      RECT 741.04 -24.64 741.36 2.2 ;
      RECT 740.77 -35.47 741.09 -25.07 ;
      RECT 739.68 -20.56 740 2.2 ;
      RECT 739 -35.52 739.32 -31.12 ;
      RECT 738.32 -35.52 738.64 2.2 ;
      RECT 737.62 -34.87 737.94 -26.325 ;
      RECT 736.96 -17.16 737.28 2.2 ;
      RECT 735.6 -17.84 735.92 2.2 ;
      RECT 735.1 -34.87 735.42 -29.475 ;
      RECT 734.24 -21.92 734.56 2.2 ;
      RECT 732.88 -18.52 733.2 2.2 ;
      RECT 732.2 -35.52 732.52 -31.12 ;
      RECT 726.08 -24.64 726.4 2.2 ;
      RECT 725.87 -35.47 726.19 -25.07 ;
      RECT 724.72 -20.56 725.04 2.2 ;
      RECT 724.04 -35.52 724.36 -31.12 ;
      RECT 723.36 -25.32 723.68 2.2 ;
      RECT 722.72 -34.87 723.04 -26.325 ;
      RECT 722 -17.16 722.32 2.2 ;
      RECT 720.64 -17.84 720.96 2.2 ;
      RECT 720.2 -34.87 720.52 -29.475 ;
      RECT 719.28 -21.92 719.6 2.2 ;
      RECT 717.92 -18.52 718.24 2.2 ;
      RECT 717.24 -35.52 717.56 -31.12 ;
      RECT 711.12 -24.64 711.44 2.2 ;
      RECT 710.97 -35.47 711.29 -25.07 ;
      RECT 709.76 -20.56 710.08 2.2 ;
      RECT 709.08 -35.52 709.4 -31.12 ;
      RECT 708.4 -25.32 708.72 2.2 ;
      RECT 707.82 -34.87 708.14 -26.325 ;
      RECT 707.04 -17.16 707.36 2.2 ;
      RECT 705.68 -17.84 706 2.2 ;
      RECT 705.3 -34.87 705.62 -29.475 ;
      RECT 704.32 -21.92 704.64 2.2 ;
      RECT 702.96 -18.52 703.28 2.2 ;
      RECT 702.28 -35.52 702.6 -31.12 ;
      RECT 696.16 -24.64 696.48 2.2 ;
      RECT 696.07 -35.47 696.39 -25.07 ;
      RECT 694.8 -20.56 695.12 2.2 ;
      RECT 694.12 -35.52 694.44 -31.12 ;
      RECT 693.44 -25.32 693.76 2.2 ;
      RECT 692.92 -34.87 693.24 -26.325 ;
      RECT 692.08 -17.16 692.4 2.2 ;
      RECT 690.72 -17.84 691.04 2.2 ;
      RECT 690.4 -34.87 690.72 -29.475 ;
      RECT 689.36 -21.92 689.68 2.2 ;
      RECT 688 -18.52 688.32 2.2 ;
      RECT 687.32 -35.52 687.64 -31.12 ;
      RECT 681.2 -20.56 681.52 2.2 ;
      RECT 681.17 -35.47 681.49 -25.07 ;
      RECT 679.84 -35.52 680.16 -31.12 ;
      RECT 679.84 -21.24 680.16 2.2 ;
      RECT 678.48 -25.32 678.8 2.2 ;
      RECT 678.02 -34.87 678.34 -26.325 ;
      RECT 677.12 -17.16 677.44 2.2 ;
      RECT 675.76 -17.84 676.08 2.2 ;
      RECT 675.5 -34.87 675.82 -29.475 ;
      RECT 674.4 -21.92 674.72 2.2 ;
      RECT 673.04 -18.52 673.36 2.2 ;
      RECT 672.36 -35.52 672.68 -31.12 ;
      RECT 666.27 -35.47 666.59 -25.07 ;
      RECT 666.24 -20.56 666.56 2.2 ;
      RECT 664.88 -35.52 665.2 -31.12 ;
      RECT 664.88 -21.24 665.2 2.2 ;
      RECT 663.52 -25.32 663.84 2.2 ;
      RECT 663.12 -34.87 663.44 -26.325 ;
      RECT 662.16 -17.16 662.48 2.2 ;
      RECT 660.8 -17.84 661.12 2.2 ;
      RECT 660.6 -34.87 660.92 -29.475 ;
      RECT 659.44 -21.92 659.76 2.2 ;
      RECT 658.08 -18.52 658.4 2.2 ;
      RECT 657.4 -35.52 657.72 -31.12 ;
      RECT 651.37 -35.47 651.69 -25.07 ;
      RECT 651.28 -20.56 651.6 2.2 ;
      RECT 649.92 -35.52 650.24 -31.12 ;
      RECT 649.92 -21.24 650.24 2.2 ;
      RECT 648.56 -25.32 648.88 2.2 ;
      RECT 648.22 -34.87 648.54 -26.325 ;
      RECT 647.2 -17.16 647.52 2.2 ;
      RECT 645.84 -17.84 646.16 2.2 ;
      RECT 645.7 -34.87 646.02 -29.475 ;
      RECT 644.48 -18.52 644.8 2.2 ;
      RECT 643.12 -21.24 643.44 2.2 ;
      RECT 642.44 -35.52 642.76 -31.12 ;
      RECT 636.47 -35.47 636.79 -25.07 ;
      RECT 636.32 -20.56 636.64 2.2 ;
      RECT 634.96 -35.52 635.28 -31.12 ;
      RECT 634.96 -21.24 635.28 2.2 ;
      RECT 633.6 -25.32 633.92 2.2 ;
      RECT 633.32 -34.87 633.64 -26.325 ;
      RECT 632.24 -17.16 632.56 2.2 ;
      RECT 630.88 -17.84 631.2 2.2 ;
      RECT 630.8 -34.87 631.12 -29.475 ;
      RECT 629.52 -18.52 629.84 2.2 ;
      RECT 628.84 -35.52 629.16 -31.12 ;
      RECT 628.16 -21.24 628.48 2.2 ;
      RECT 621.57 -35.47 621.89 -25.07 ;
      RECT 621.36 -20.56 621.68 2.2 ;
      RECT 620 -35.52 620.32 -31.12 ;
      RECT 620 -21.24 620.32 2.2 ;
      RECT 618.64 -25.32 618.96 2.2 ;
      RECT 618.42 -34.87 618.74 -26.325 ;
      RECT 617.28 -17.16 617.6 2.2 ;
      RECT 615.92 -17.84 616.24 2.2 ;
      RECT 615.9 -34.87 616.22 -29.475 ;
      RECT 614.56 -18.52 614.88 2.2 ;
      RECT 613.88 -35.52 614.2 -31.12 ;
      RECT 613.2 -21.24 613.52 2.2 ;
      RECT 606.67 -35.47 606.99 -25.07 ;
      RECT 606.4 -20.56 606.72 2.2 ;
      RECT 605.04 -35.52 605.36 -31.12 ;
      RECT 605.04 -21.24 605.36 2.2 ;
      RECT 603.68 -25.32 604 2.2 ;
      RECT 603.52 -34.87 603.84 -26.325 ;
      RECT 602.32 -17.16 602.64 2.2 ;
      RECT 601 -34.87 601.32 -29.475 ;
      RECT 600.96 -17.84 601.28 2.2 ;
      RECT 599.6 -18.52 599.92 2.2 ;
      RECT 598.92 -35.52 599.24 -31.12 ;
      RECT 598.24 -21.24 598.56 2.2 ;
      RECT 591.77 -35.47 592.09 -25.07 ;
      RECT 591.44 -20.56 591.76 2.2 ;
      RECT 590.08 -35.52 590.4 -31.12 ;
      RECT 590.08 -21.24 590.4 2.2 ;
      RECT 588.72 -25.32 589.04 2.2 ;
      RECT 588.62 -34.87 588.94 -26.325 ;
      RECT 587.36 -17.16 587.68 2.2 ;
      RECT 586.1 -34.87 586.42 -29.475 ;
      RECT 586 -18.52 586.32 2.2 ;
      RECT 584.64 -18.52 584.96 2.2 ;
      RECT 583.96 -35.52 584.28 -31.12 ;
      RECT 583.28 -21.24 583.6 2.2 ;
      RECT 576.87 -35.47 577.19 -25.07 ;
      RECT 576.48 -20.56 576.8 2.2 ;
      RECT 575.12 -35.52 575.44 -31.12 ;
      RECT 575.12 -21.24 575.44 2.2 ;
      RECT 573.76 -25.32 574.08 2.2 ;
      RECT 573.72 -34.87 574.04 -26.325 ;
      RECT 572.4 -17.16 572.72 2.2 ;
      RECT 571.2 -34.87 571.52 -29.475 ;
      RECT 571.04 -18.52 571.36 2.2 ;
      RECT 569.68 -18.52 570 2.2 ;
      RECT 569 -35.52 569.32 -31.12 ;
      RECT 568.32 -21.24 568.64 2.2 ;
      RECT 561.97 -35.47 562.29 -25.07 ;
      RECT 561.52 -20.56 561.84 2.2 ;
      RECT 560.16 -35.52 560.48 -31.12 ;
      RECT 560.16 -21.24 560.48 2.2 ;
      RECT 558.82 -34.87 559.14 -26.325 ;
      RECT 558.8 -25.32 559.12 2.2 ;
      RECT 557.44 -17.16 557.76 2.2 ;
      RECT 556.3 -34.87 556.62 -29.475 ;
      RECT 556.08 -18.52 556.4 2.2 ;
      RECT 554.72 -18.52 555.04 2.2 ;
      RECT 554.04 -35.52 554.36 -31.12 ;
      RECT 553.36 -21.24 553.68 2.2 ;
      RECT 547.07 -35.47 547.39 -25.07 ;
      RECT 546.56 -20.56 546.88 2.2 ;
      RECT 545.2 -35.52 545.52 -31.12 ;
      RECT 545.2 -21.24 545.52 2.2 ;
      RECT 543.92 -34.87 544.24 -26.325 ;
      RECT 543.84 -25.32 544.16 2.2 ;
      RECT 542.48 -17.16 542.8 2.2 ;
      RECT 541.4 -34.87 541.72 -29.475 ;
      RECT 541.12 -18.52 541.44 2.2 ;
      RECT 539.76 -18.52 540.08 2.2 ;
      RECT 539.08 -35.52 539.4 -31.12 ;
      RECT 538.4 -21.24 538.72 2.2 ;
      RECT 532.17 -35.47 532.49 -25.07 ;
      RECT 531.6 -20.56 531.92 2.2 ;
      RECT 530.24 -35.52 530.56 -31.12 ;
      RECT 530.24 -21.24 530.56 2.2 ;
      RECT 529.02 -34.87 529.34 -26.325 ;
      RECT 528.88 -25.32 529.2 2.2 ;
      RECT 527.52 -17.16 527.84 2.2 ;
      RECT 526.5 -34.87 526.82 -29.475 ;
      RECT 526.16 -18.52 526.48 2.2 ;
      RECT 524.8 -18.52 525.12 2.2 ;
      RECT 524.12 -35.52 524.44 -31.12 ;
      RECT 523.44 -21.24 523.76 2.2 ;
      RECT 517.27 -35.47 517.59 -25.07 ;
      RECT 516.64 -20.56 516.96 2.2 ;
      RECT 515.96 -35.52 516.28 -31.12 ;
      RECT 515.28 -35.52 515.6 2.2 ;
      RECT 514.12 -34.87 514.44 -26.325 ;
      RECT 513.92 -25.32 514.24 2.2 ;
      RECT 512.56 -17.16 512.88 2.2 ;
      RECT 511.6 -34.87 511.92 -29.475 ;
      RECT 511.2 -18.52 511.52 2.2 ;
      RECT 509.84 -18.52 510.16 2.2 ;
      RECT 509.16 -35.52 509.48 -31.12 ;
      RECT 508.48 -21.24 508.8 2.2 ;
      RECT 503.04 -24.64 503.36 2.2 ;
      RECT 502.37 -35.47 502.69 -25.07 ;
      RECT 501.68 -20.56 502 2.2 ;
      RECT 501 -35.52 501.32 -31.12 ;
      RECT 500.32 -35.52 500.64 2.2 ;
      RECT 499.22 -34.87 499.54 -26.325 ;
      RECT 498.96 -25.32 499.28 2.2 ;
      RECT 497.6 -17.16 497.92 2.2 ;
      RECT 496.7 -34.87 497.02 -29.475 ;
      RECT 496.24 -18.52 496.56 2.2 ;
      RECT 494.88 -18.52 495.2 2.2 ;
      RECT 494.2 -35.52 494.52 -31.12 ;
      RECT 493.52 -21.24 493.84 2.2 ;
      RECT 488.08 -24.64 488.4 2.2 ;
      RECT 487.47 -35.47 487.79 -25.07 ;
      RECT 486.72 -20.56 487.04 2.2 ;
      RECT 486.04 -35.52 486.36 -31.12 ;
      RECT 485.36 -35.52 485.68 2.2 ;
      RECT 484.32 -34.87 484.64 -26.325 ;
      RECT 484 -25.32 484.32 2.2 ;
      RECT 482.64 -17.16 482.96 2.2 ;
      RECT 481.8 -34.87 482.12 -29.475 ;
      RECT 481.28 -18.52 481.6 2.2 ;
      RECT 479.92 -18.52 480.24 2.2 ;
      RECT 479.24 -35.52 479.56 -31.12 ;
      RECT 478.56 -21.24 478.88 2.2 ;
      RECT 473.12 -24.64 473.44 2.2 ;
      RECT 472.57 -35.47 472.89 -25.07 ;
      RECT 471.76 -20.56 472.08 2.2 ;
      RECT 471.08 -35.52 471.4 -31.12 ;
      RECT 470.4 -35.52 470.72 2.2 ;
      RECT 469.42 -34.87 469.74 -26.325 ;
      RECT 469.04 -25.32 469.36 2.2 ;
      RECT 467.68 -17.16 468 2.2 ;
      RECT 466.9 -34.87 467.22 -29.475 ;
      RECT 466.32 -18.52 466.64 2.2 ;
      RECT 464.96 -35.52 465.28 -30.44 ;
      RECT 464.96 -18.52 465.28 2.2 ;
      RECT 464.28 -35.52 464.6 -31.12 ;
      RECT 458.16 -24.64 458.48 2.2 ;
      RECT 457.67 -35.47 457.99 -25.07 ;
      RECT 456.8 -20.56 457.12 2.2 ;
      RECT 456.12 -35.52 456.44 -31.12 ;
      RECT 455.44 -35.52 455.76 2.2 ;
      RECT 454.52 -34.87 454.84 -26.325 ;
      RECT 454.08 -25.32 454.4 2.2 ;
      RECT 452.72 -17.16 453.04 2.2 ;
      RECT 452 -34.87 452.32 -29.475 ;
      RECT 451.36 -18.52 451.68 2.2 ;
      RECT 450 -18.52 450.32 2.2 ;
      RECT 449.32 -35.52 449.64 -31.12 ;
      RECT 443.2 -24.64 443.52 2.2 ;
      RECT 442.77 -35.47 443.09 -25.07 ;
      RECT 441.84 -20.56 442.16 2.2 ;
      RECT 441.16 -35.52 441.48 -31.12 ;
      RECT 440.48 -35.52 440.8 2.2 ;
      RECT 439.62 -34.87 439.94 -26.325 ;
      RECT 439.12 -25.32 439.44 2.2 ;
      RECT 437.76 -17.16 438.08 2.2 ;
      RECT 437.1 -34.87 437.42 -29.475 ;
      RECT 436.4 -21.92 436.72 2.2 ;
      RECT 435.04 -18.52 435.36 2.2 ;
      RECT 434.36 -35.52 434.68 -31.12 ;
      RECT 428.24 -24.64 428.56 2.2 ;
      RECT 427.87 -35.47 428.19 -25.07 ;
      RECT 426.88 -20.56 427.2 2.2 ;
      RECT 426.2 -35.52 426.52 -31.12 ;
      RECT 425.52 -35.52 425.84 2.2 ;
      RECT 424.72 -34.87 425.04 -26.325 ;
      RECT 424.16 -25.32 424.48 2.2 ;
      RECT 422.8 -17.16 423.12 2.2 ;
      RECT 422.2 -34.87 422.52 -29.475 ;
      RECT 421.44 -21.92 421.76 2.2 ;
      RECT 420.08 -18.52 420.4 2.2 ;
      RECT 419.4 -35.52 419.72 -31.12 ;
      RECT 413.28 -24.64 413.6 2.2 ;
      RECT 412.97 -35.47 413.29 -25.07 ;
      RECT 411.92 -20.56 412.24 2.2 ;
      RECT 411.24 -35.52 411.56 -31.12 ;
      RECT 410.56 -35.52 410.88 2.2 ;
      RECT 409.82 -34.87 410.14 -26.325 ;
      RECT 409.2 -17.16 409.52 2.2 ;
      RECT 407.84 -17.84 408.16 2.2 ;
      RECT 407.3 -34.87 407.62 -29.475 ;
      RECT 406.48 -21.92 406.8 2.2 ;
      RECT 405.12 -18.52 405.44 2.2 ;
      RECT 404.44 -35.52 404.76 -31.12 ;
      RECT 398.32 -24.64 398.64 2.2 ;
      RECT 398.07 -35.47 398.39 -25.07 ;
      RECT 396.96 -20.56 397.28 2.2 ;
      RECT 396.28 -35.52 396.6 -31.12 ;
      RECT 395.6 -35.52 395.92 2.2 ;
      RECT 394.92 -34.87 395.24 -26.325 ;
      RECT 394.24 -17.16 394.56 2.2 ;
      RECT 392.88 -17.84 393.2 2.2 ;
      RECT 392.4 -34.87 392.72 -29.475 ;
      RECT 391.52 -21.92 391.84 2.2 ;
      RECT 390.16 -18.52 390.48 2.2 ;
      RECT 389.48 -35.52 389.8 -31.12 ;
      RECT 383.36 -24.64 383.68 2.2 ;
      RECT 383.17 -35.47 383.49 -25.07 ;
      RECT 382 -20.56 382.32 2.2 ;
      RECT 381.32 -35.52 381.64 -31.12 ;
      RECT 380.64 -25.32 380.96 2.2 ;
      RECT 380.02 -34.87 380.34 -26.325 ;
      RECT 379.28 -17.16 379.6 2.2 ;
      RECT 377.92 -17.84 378.24 2.2 ;
      RECT 377.5 -34.87 377.82 -29.475 ;
      RECT 376.56 -21.92 376.88 2.2 ;
      RECT 375.2 -18.52 375.52 2.2 ;
      RECT 374.52 -35.52 374.84 -31.12 ;
      RECT 368.4 -24.64 368.72 2.2 ;
      RECT 368.27 -35.47 368.59 -25.07 ;
      RECT 367.04 -20.56 367.36 2.2 ;
      RECT 366.36 -35.52 366.68 -31.12 ;
      RECT 365.68 -25.32 366 2.2 ;
      RECT 365.12 -34.87 365.44 -26.325 ;
      RECT 364.32 -17.16 364.64 2.2 ;
      RECT 362.96 -17.84 363.28 2.2 ;
      RECT 362.6 -34.87 362.92 -29.475 ;
      RECT 361.6 -21.92 361.92 2.2 ;
      RECT 360.24 -18.52 360.56 2.2 ;
      RECT 359.56 -35.52 359.88 -31.12 ;
      RECT 353.44 -24.64 353.76 2.2 ;
      RECT 353.37 -35.47 353.69 -25.07 ;
      RECT 352.08 -20.56 352.4 2.2 ;
      RECT 350.72 -25.32 351.04 2.2 ;
      RECT 350.22 -34.87 350.54 -26.325 ;
      RECT 349.36 -17.16 349.68 2.2 ;
      RECT 348 -17.84 348.32 2.2 ;
      RECT 347.7 -34.87 348.02 -29.475 ;
      RECT 346.64 -21.92 346.96 2.2 ;
      RECT 345.28 -18.52 345.6 2.2 ;
      RECT 344.6 -35.52 344.92 -31.12 ;
      RECT 338.48 -20.56 338.8 2.2 ;
      RECT 338.47 -35.47 338.79 -25.07 ;
      RECT 337.12 -35.52 337.44 -31.12 ;
      RECT 337.12 -21.24 337.44 2.2 ;
      RECT 335.76 -25.32 336.08 2.2 ;
      RECT 335.32 -34.87 335.64 -26.325 ;
      RECT 334.4 -17.16 334.72 2.2 ;
      RECT 333.04 -17.84 333.36 2.2 ;
      RECT 332.8 -34.87 333.12 -29.475 ;
      RECT 331.68 -21.92 332 2.2 ;
      RECT 330.32 -18.52 330.64 2.2 ;
      RECT 329.64 -35.52 329.96 -31.12 ;
      RECT 323.57 -35.47 323.89 -25.07 ;
      RECT 323.52 -20.56 323.84 2.2 ;
      RECT 322.16 -35.52 322.48 -31.12 ;
      RECT 322.16 -21.24 322.48 2.2 ;
      RECT 320.8 -25.32 321.12 2.2 ;
      RECT 320.42 -34.87 320.74 -26.325 ;
      RECT 319.44 -17.16 319.76 2.2 ;
      RECT 318.08 -17.84 318.4 2.2 ;
      RECT 317.9 -34.87 318.22 -29.475 ;
      RECT 316.72 -21.92 317.04 2.2 ;
      RECT 315.36 -18.52 315.68 2.2 ;
      RECT 314.68 -35.52 315 -31.12 ;
      RECT 308.67 -35.47 308.99 -25.07 ;
      RECT 308.56 -20.56 308.88 2.2 ;
      RECT 307.2 -35.52 307.52 -31.12 ;
      RECT 307.2 -21.24 307.52 2.2 ;
      RECT 305.84 -25.32 306.16 2.2 ;
      RECT 305.52 -34.87 305.84 -26.325 ;
      RECT 304.48 -17.16 304.8 2.2 ;
      RECT 303.12 -17.84 303.44 2.2 ;
      RECT 303 -34.87 303.32 -29.475 ;
      RECT 301.76 -18.52 302.08 2.2 ;
      RECT 300.4 -21.24 300.72 2.2 ;
      RECT 299.72 -35.52 300.04 -31.12 ;
      RECT 293.77 -35.47 294.09 -25.07 ;
      RECT 293.6 -20.56 293.92 2.2 ;
      RECT 292.24 -35.52 292.56 -31.12 ;
      RECT 292.24 -21.24 292.56 2.2 ;
      RECT 290.88 -25.32 291.2 2.2 ;
      RECT 290.62 -34.87 290.94 -26.325 ;
      RECT 289.52 -17.16 289.84 2.2 ;
      RECT 288.16 -17.84 288.48 2.2 ;
      RECT 288.1 -34.87 288.42 -29.475 ;
      RECT 286.8 -18.52 287.12 2.2 ;
      RECT 286.12 -35.52 286.44 -31.12 ;
      RECT 285.44 -21.24 285.76 2.2 ;
      RECT 278.87 -35.47 279.19 -25.07 ;
      RECT 278.64 -20.56 278.96 2.2 ;
      RECT 277.28 -35.52 277.6 -31.12 ;
      RECT 277.28 -21.24 277.6 2.2 ;
      RECT 275.92 -25.32 276.24 2.2 ;
      RECT 275.72 -34.87 276.04 -26.325 ;
      RECT 274.56 -17.16 274.88 2.2 ;
      RECT 273.2 -34.87 273.52 -29.475 ;
      RECT 273.2 -17.84 273.52 2.2 ;
      RECT 271.84 -18.52 272.16 2.2 ;
      RECT 271.16 -35.52 271.48 -31.12 ;
      RECT 270.48 -21.24 270.8 2.2 ;
      RECT 263.97 -35.47 264.29 -25.07 ;
      RECT 263.68 -20.56 264 2.2 ;
      RECT 262.32 -35.52 262.64 -31.12 ;
      RECT 262.32 -21.24 262.64 2.2 ;
      RECT 260.96 -25.32 261.28 2.2 ;
      RECT 260.82 -34.87 261.14 -26.325 ;
      RECT 259.6 -17.16 259.92 2.2 ;
      RECT 258.3 -34.87 258.62 -29.475 ;
      RECT 258.24 -18.52 258.56 2.2 ;
      RECT 256.88 -18.52 257.2 2.2 ;
      RECT 256.2 -35.52 256.52 -31.12 ;
      RECT 255.52 -21.24 255.84 2.2 ;
      RECT 249.07 -35.47 249.39 -25.07 ;
      RECT 248.72 -20.56 249.04 2.2 ;
      RECT 247.36 -35.52 247.68 -31.12 ;
      RECT 247.36 -21.24 247.68 2.2 ;
      RECT 246 -25.32 246.32 2.2 ;
      RECT 245.92 -34.87 246.24 -26.325 ;
      RECT 244.64 -17.16 244.96 2.2 ;
      RECT 243.4 -34.87 243.72 -29.475 ;
      RECT 243.28 -18.52 243.6 2.2 ;
      RECT 241.92 -18.52 242.24 2.2 ;
      RECT 241.24 -35.52 241.56 -31.12 ;
      RECT 240.56 -21.24 240.88 2.2 ;
      RECT 234.17 -35.47 234.49 -25.07 ;
      RECT 233.76 -20.56 234.08 2.2 ;
      RECT 232.4 -35.52 232.72 -31.12 ;
      RECT 232.4 -21.24 232.72 2.2 ;
      RECT 231.04 -25.32 231.36 2.2 ;
      RECT 231.02 -34.87 231.34 -26.325 ;
      RECT 229.68 -17.16 230 2.2 ;
      RECT 228.5 -34.87 228.82 -29.475 ;
      RECT 228.32 -18.52 228.64 2.2 ;
      RECT 226.96 -18.52 227.28 2.2 ;
      RECT 226.28 -35.52 226.6 -31.12 ;
      RECT 225.6 -21.24 225.92 2.2 ;
      RECT 219.27 -35.47 219.59 -25.07 ;
      RECT 218.8 -20.56 219.12 2.2 ;
      RECT 217.44 -35.52 217.76 -31.12 ;
      RECT 217.44 -21.24 217.76 2.2 ;
      RECT 216.12 -34.87 216.44 -26.325 ;
      RECT 216.08 -25.32 216.4 2.2 ;
      RECT 214.72 -17.16 215.04 2.2 ;
      RECT 213.6 -34.87 213.92 -29.475 ;
      RECT 213.36 -18.52 213.68 2.2 ;
      RECT 212 -18.52 212.32 2.2 ;
      RECT 211.32 -35.52 211.64 -31.12 ;
      RECT 210.64 -21.24 210.96 2.2 ;
      RECT 204.37 -35.47 204.69 -25.07 ;
      RECT 203.84 -20.56 204.16 2.2 ;
      RECT 202.48 -35.52 202.8 -31.12 ;
      RECT 202.48 -21.24 202.8 2.2 ;
      RECT 201.22 -34.87 201.54 -26.325 ;
      RECT 201.12 -25.32 201.44 2.2 ;
      RECT 199.76 -17.16 200.08 2.2 ;
      RECT 198.7 -34.87 199.02 -29.475 ;
      RECT 198.4 -18.52 198.72 2.2 ;
      RECT 197.04 -18.52 197.36 2.2 ;
      RECT 196.36 -35.52 196.68 -31.12 ;
      RECT 195.68 -21.24 196 2.2 ;
      RECT 189.47 -35.47 189.79 -25.07 ;
      RECT 188.88 -20.56 189.2 2.2 ;
      RECT 187.52 -35.52 187.84 -31.12 ;
      RECT 187.52 -21.24 187.84 2.2 ;
      RECT 186.32 -34.87 186.64 -26.325 ;
      RECT 186.16 -25.32 186.48 2.2 ;
      RECT 184.8 -17.16 185.12 2.2 ;
      RECT 183.8 -34.87 184.12 -29.475 ;
      RECT 183.44 -18.52 183.76 2.2 ;
      RECT 182.08 -18.52 182.4 2.2 ;
      RECT 181.4 -35.52 181.72 -31.12 ;
      RECT 180.72 -21.24 181.04 2.2 ;
      RECT 174.57 -35.47 174.89 -25.07 ;
      RECT 173.92 -20.56 174.24 2.2 ;
      RECT 173.24 -35.52 173.56 -31.12 ;
      RECT 172.56 -35.52 172.88 2.2 ;
      RECT 171.42 -34.87 171.74 -26.325 ;
      RECT 171.2 -25.32 171.52 2.2 ;
      RECT 169.84 -17.16 170.16 2.2 ;
      RECT 168.9 -34.87 169.22 -29.475 ;
      RECT 168.48 -18.52 168.8 2.2 ;
      RECT 167.12 -18.52 167.44 2.2 ;
      RECT 166.44 -35.52 166.76 -31.12 ;
      RECT 165.76 -21.24 166.08 2.2 ;
      RECT 160.32 -24.64 160.64 2.2 ;
      RECT 159.67 -35.47 159.99 -25.07 ;
      RECT 158.96 -20.56 159.28 2.2 ;
      RECT 158.28 -35.52 158.6 -31.12 ;
      RECT 157.6 -35.52 157.92 2.2 ;
      RECT 156.52 -34.87 156.84 -26.325 ;
      RECT 156.24 -25.32 156.56 2.2 ;
      RECT 154.88 -17.16 155.2 2.2 ;
      RECT 154 -34.87 154.32 -29.475 ;
      RECT 153.52 -18.52 153.84 2.2 ;
      RECT 152.16 -18.52 152.48 2.2 ;
      RECT 151.48 -35.52 151.8 -31.12 ;
      RECT 150.8 -21.24 151.12 2.2 ;
      RECT 145.36 -24.64 145.68 2.2 ;
      RECT 144.77 -35.47 145.09 -25.07 ;
      RECT 144 -20.56 144.32 2.2 ;
      RECT 143.32 -35.52 143.64 -31.12 ;
      RECT 142.64 -35.52 142.96 2.2 ;
      RECT 141.62 -34.87 141.94 -26.325 ;
      RECT 141.28 -25.32 141.6 2.2 ;
      RECT 139.92 -17.16 140.24 2.2 ;
      RECT 139.1 -34.87 139.42 -29.475 ;
      RECT 138.56 -18.52 138.88 2.2 ;
      RECT 137.2 -18.52 137.52 2.2 ;
      RECT 136.52 -35.52 136.84 -31.12 ;
      RECT 135.84 -21.24 136.16 2.2 ;
      RECT 130.4 -24.64 130.72 2.2 ;
      RECT 129.87 -35.47 130.19 -25.07 ;
      RECT 129.04 -20.56 129.36 2.2 ;
      RECT 128.36 -35.52 128.68 -31.12 ;
      RECT 127.68 -35.52 128 2.2 ;
      RECT 126.72 -34.87 127.04 -26.325 ;
      RECT 126.32 -25.32 126.64 2.2 ;
      RECT 124.96 -17.16 125.28 2.2 ;
      RECT 124.2 -34.87 124.52 -29.475 ;
      RECT 123.6 -18.52 123.92 2.2 ;
      RECT 122.24 -18.52 122.56 2.2 ;
      RECT 121.56 -35.52 121.88 -31.12 ;
      RECT 115.44 -24.64 115.76 2.2 ;
      RECT 114.97 -35.47 115.29 -25.07 ;
      RECT 114.08 -20.56 114.4 2.2 ;
      RECT 113.4 -35.52 113.72 -31.12 ;
      RECT 112.72 -35.52 113.04 2.2 ;
      RECT 111.82 -34.87 112.14 -26.325 ;
      RECT 111.36 -25.32 111.68 2.2 ;
      RECT 110 -17.16 110.32 2.2 ;
      RECT 109.3 -34.87 109.62 -29.475 ;
      RECT 108.64 -18.52 108.96 2.2 ;
      RECT 107.28 -18.52 107.6 2.2 ;
      RECT 106.6 -35.52 106.92 -31.12 ;
      RECT 100.48 -24.64 100.8 2.2 ;
      RECT 100.07 -35.47 100.39 -25.07 ;
      RECT 99.12 -20.56 99.44 2.2 ;
      RECT 98.44 -35.52 98.76 -31.12 ;
      RECT 97.76 -35.52 98.08 2.2 ;
      RECT 96.92 -34.87 97.24 -26.325 ;
      RECT 96.4 -25.32 96.72 2.2 ;
      RECT 95.04 -17.16 95.36 2.2 ;
      RECT 94.4 -34.87 94.72 -29.475 ;
      RECT 93.68 -21.92 94 2.2 ;
      RECT 92.32 -18.52 92.64 2.2 ;
      RECT 91.64 -35.52 91.96 -31.12 ;
      RECT 85.52 -24.64 85.84 2.2 ;
      RECT 85.17 -35.47 85.49 -25.07 ;
      RECT 84.16 -20.56 84.48 2.2 ;
      RECT 83.48 -35.52 83.8 -31.12 ;
      RECT 82.8 -35.52 83.12 2.2 ;
      RECT 82.02 -34.87 82.34 -26.325 ;
      RECT 81.44 -25.32 81.76 2.2 ;
      RECT 80.08 -17.84 80.4 2.2 ;
      RECT 79.5 -34.87 79.82 -29.475 ;
      RECT 78.72 -21.92 79.04 2.2 ;
      RECT 77.36 -18.52 77.68 2.2 ;
      RECT 76.68 -35.52 77 -31.12 ;
      RECT 70.56 -24.64 70.88 2.2 ;
      RECT 70.27 -35.47 70.59 -25.07 ;
      RECT 69.2 -20.56 69.52 2.2 ;
      RECT 68.52 -35.52 68.84 -31.12 ;
      RECT 67.84 -35.52 68.16 2.2 ;
      RECT 67.12 -34.87 67.44 -26.325 ;
      RECT 66.48 -17.16 66.8 2.2 ;
      RECT 65.12 -17.84 65.44 2.2 ;
      RECT 64.6 -34.87 64.92 -29.475 ;
      RECT 63.76 -21.92 64.08 2.2 ;
      RECT 62.4 -18.52 62.72 2.2 ;
      RECT 61.72 -35.52 62.04 -31.12 ;
      RECT 55.6 -24.64 55.92 2.2 ;
      RECT 55.37 -35.47 55.69 -25.07 ;
      RECT 54.24 -20.56 54.56 2.2 ;
      RECT 53.56 -35.52 53.88 -31.12 ;
      RECT 52.88 -25.32 53.2 2.2 ;
      RECT 52.22 -34.87 52.54 -26.325 ;
      RECT 51.52 -17.16 51.84 2.2 ;
      RECT 50.16 -17.84 50.48 2.2 ;
      RECT 49.7 -34.87 50.02 -29.475 ;
      RECT 48.8 -21.92 49.12 2.2 ;
      RECT 47.44 -18.52 47.76 2.2 ;
      RECT 46.76 -35.52 47.08 -31.12 ;
      RECT 40.64 -24.64 40.96 2.2 ;
      RECT 40.47 -35.47 40.79 -25.07 ;
      RECT 39.28 -20.56 39.6 2.2 ;
      RECT 38.6 -35.52 38.92 -31.12 ;
      RECT 37.92 -25.32 38.24 2.2 ;
      RECT 37.32 -34.87 37.64 -26.325 ;
      RECT 36.56 -17.16 36.88 2.2 ;
      RECT 35.2 -17.84 35.52 2.2 ;
      RECT 34.8 -34.87 35.12 -29.475 ;
      RECT 33.84 -21.92 34.16 2.2 ;
      RECT 32.48 -18.52 32.8 2.2 ;
      RECT 31.8 -35.52 32.12 -31.12 ;
      RECT 25.68 -24.64 26 2.2 ;
      RECT 25.57 -35.47 25.89 -25.07 ;
      RECT 24.32 -20.56 24.64 2.2 ;
      RECT 23.64 -35.52 23.96 -31.12 ;
      RECT 22.96 -25.32 23.28 2.2 ;
      RECT 22.42 -34.87 22.74 -26.325 ;
      RECT 21.6 -17.16 21.92 2.2 ;
      RECT 20.24 -17.84 20.56 2.2 ;
      RECT 19.9 -34.87 20.22 -29.475 ;
      RECT 18.88 -21.92 19.2 2.2 ;
      RECT 17.52 -18.52 17.84 2.2 ;
      RECT 16.84 -35.52 17.16 -31.12 ;
      RECT 10.04 -35.47 10.36 -21.29 ;
      RECT 9.36 -21.24 9.68 2.2 ;
      RECT 8 -34.16 8.32 2.2 ;
      RECT 6.64 -34.16 6.96 2.2 ;
      RECT 5.28 -17.84 5.6 2.2 ;
      RECT 4.6 -35.52 4.92 -23.64 ;
      RECT 3.92 -21.92 4.24 2.2 ;
      RECT 3.24 -35.52 3.56 -25 ;
      RECT 2.56 -21.24 2.88 2.2 ;
      RECT 1.88 -35.52 2.2 -25.68 ;
    LAYER met2 SPACING 0.14 ;
      RECT -1.525 -34.8 954.885 2.225 ;
      RECT 946.865 -35.545 954.885 2.225 ;
      RECT 945.585 -34.82 954.885 2.225 ;
      RECT 945.605 -34.825 954.885 2.225 ;
      RECT 928.165 -34.82 944.655 2.225 ;
      RECT 913.265 -34.82 927.235 2.225 ;
      RECT 898.365 -34.82 912.335 2.225 ;
      RECT 883.465 -34.82 897.435 2.225 ;
      RECT 868.565 -34.82 882.535 2.225 ;
      RECT 853.665 -34.82 867.635 2.225 ;
      RECT 838.765 -34.82 852.735 2.225 ;
      RECT 823.865 -34.82 837.835 2.225 ;
      RECT 808.965 -34.82 822.935 2.225 ;
      RECT 794.065 -34.82 808.035 2.225 ;
      RECT 779.165 -34.82 793.135 2.225 ;
      RECT 764.265 -34.82 778.235 2.225 ;
      RECT 749.365 -34.82 763.335 2.225 ;
      RECT 734.465 -34.82 748.435 2.225 ;
      RECT 719.565 -34.82 733.535 2.225 ;
      RECT 704.665 -34.82 718.635 2.225 ;
      RECT 689.765 -34.82 703.735 2.225 ;
      RECT 674.865 -34.82 688.835 2.225 ;
      RECT 659.965 -34.82 673.935 2.225 ;
      RECT 645.065 -34.82 659.035 2.225 ;
      RECT 630.165 -34.82 644.135 2.225 ;
      RECT 615.265 -34.82 629.235 2.225 ;
      RECT 600.365 -34.82 614.335 2.225 ;
      RECT 585.465 -34.82 599.435 2.225 ;
      RECT 570.565 -34.82 584.535 2.225 ;
      RECT 555.665 -34.82 569.635 2.225 ;
      RECT 540.765 -34.82 554.735 2.225 ;
      RECT 525.865 -34.82 539.835 2.225 ;
      RECT 510.965 -34.82 524.935 2.225 ;
      RECT 496.065 -34.82 510.035 2.225 ;
      RECT 481.165 -34.82 495.135 2.225 ;
      RECT 466.265 -34.82 480.235 2.225 ;
      RECT 451.365 -34.82 465.335 2.225 ;
      RECT 436.465 -34.82 450.435 2.225 ;
      RECT 421.565 -34.82 435.535 2.225 ;
      RECT 406.665 -34.82 420.635 2.225 ;
      RECT 391.765 -34.82 405.735 2.225 ;
      RECT 376.865 -34.82 390.835 2.225 ;
      RECT 361.965 -34.82 375.935 2.225 ;
      RECT 347.065 -34.82 361.035 2.225 ;
      RECT 332.165 -34.82 346.135 2.225 ;
      RECT 317.265 -34.82 331.235 2.225 ;
      RECT 302.365 -34.82 316.335 2.225 ;
      RECT 287.465 -34.82 301.435 2.225 ;
      RECT 272.565 -34.82 286.535 2.225 ;
      RECT 257.665 -34.82 271.635 2.225 ;
      RECT 242.765 -34.82 256.735 2.225 ;
      RECT 227.865 -34.82 241.835 2.225 ;
      RECT 212.965 -34.82 226.935 2.225 ;
      RECT 198.065 -34.82 212.035 2.225 ;
      RECT 183.165 -34.82 197.135 2.225 ;
      RECT 168.265 -34.82 182.235 2.225 ;
      RECT 153.365 -34.82 167.335 2.225 ;
      RECT 138.465 -34.82 152.435 2.225 ;
      RECT 123.565 -34.82 137.535 2.225 ;
      RECT 108.665 -34.82 122.635 2.225 ;
      RECT 93.765 -34.82 107.735 2.225 ;
      RECT 78.865 -34.82 92.835 2.225 ;
      RECT 63.965 -34.82 77.935 2.225 ;
      RECT 49.065 -34.82 63.035 2.225 ;
      RECT 34.165 -34.82 48.135 2.225 ;
      RECT 19.265 -34.82 33.235 2.225 ;
      RECT 6.885 -34.82 18.335 2.225 ;
      RECT -1.525 -34.82 5.955 2.225 ;
      RECT 928.185 -34.825 944.635 2.225 ;
      RECT 931.965 -35.545 944.635 2.225 ;
      RECT 913.285 -34.825 927.215 2.225 ;
      RECT 917.065 -35.545 927.215 2.225 ;
      RECT 898.385 -34.825 912.315 2.225 ;
      RECT 902.165 -35.545 912.315 2.225 ;
      RECT 883.485 -34.825 897.415 2.225 ;
      RECT 887.265 -35.545 897.415 2.225 ;
      RECT 868.585 -34.825 882.515 2.225 ;
      RECT 872.365 -35.545 882.515 2.225 ;
      RECT 853.685 -34.825 867.615 2.225 ;
      RECT 857.465 -35.545 867.615 2.225 ;
      RECT 838.785 -34.825 852.715 2.225 ;
      RECT 842.565 -35.545 852.715 2.225 ;
      RECT 823.885 -34.825 837.815 2.225 ;
      RECT 827.665 -35.545 837.815 2.225 ;
      RECT 808.985 -34.825 822.915 2.225 ;
      RECT 812.765 -35.545 822.915 2.225 ;
      RECT 794.085 -34.825 808.015 2.225 ;
      RECT 797.865 -35.545 808.015 2.225 ;
      RECT 779.185 -34.825 793.115 2.225 ;
      RECT 782.965 -35.545 793.115 2.225 ;
      RECT 764.285 -34.825 778.215 2.225 ;
      RECT 768.065 -35.545 778.215 2.225 ;
      RECT 749.385 -34.825 763.315 2.225 ;
      RECT 753.165 -35.545 763.315 2.225 ;
      RECT 734.485 -34.825 748.415 2.225 ;
      RECT 738.265 -35.545 748.415 2.225 ;
      RECT 719.585 -34.825 733.515 2.225 ;
      RECT 723.365 -35.545 733.515 2.225 ;
      RECT 704.685 -34.825 718.615 2.225 ;
      RECT 708.465 -35.545 718.615 2.225 ;
      RECT 689.785 -34.825 703.715 2.225 ;
      RECT 693.565 -35.545 703.715 2.225 ;
      RECT 674.885 -34.825 688.815 2.225 ;
      RECT 678.665 -35.545 688.815 2.225 ;
      RECT 659.985 -34.825 673.915 2.225 ;
      RECT 663.765 -35.545 673.915 2.225 ;
      RECT 645.085 -34.825 659.015 2.225 ;
      RECT 648.865 -35.545 659.015 2.225 ;
      RECT 630.185 -34.825 644.115 2.225 ;
      RECT 633.965 -35.545 644.115 2.225 ;
      RECT 615.285 -34.825 629.215 2.225 ;
      RECT 619.065 -35.545 629.215 2.225 ;
      RECT 600.385 -34.825 614.315 2.225 ;
      RECT 604.165 -35.545 614.315 2.225 ;
      RECT 585.485 -34.825 599.415 2.225 ;
      RECT 589.265 -35.545 599.415 2.225 ;
      RECT 570.585 -34.825 584.515 2.225 ;
      RECT 574.365 -35.545 584.515 2.225 ;
      RECT 555.685 -34.825 569.615 2.225 ;
      RECT 559.465 -35.545 569.615 2.225 ;
      RECT 540.785 -34.825 554.715 2.225 ;
      RECT 544.565 -35.545 554.715 2.225 ;
      RECT 525.885 -34.825 539.815 2.225 ;
      RECT 529.665 -35.545 539.815 2.225 ;
      RECT 510.985 -34.825 524.915 2.225 ;
      RECT 514.765 -35.545 524.915 2.225 ;
      RECT 496.085 -34.825 510.015 2.225 ;
      RECT 499.865 -35.545 510.015 2.225 ;
      RECT 481.185 -34.825 495.115 2.225 ;
      RECT 484.965 -35.545 495.115 2.225 ;
      RECT 466.285 -34.825 480.215 2.225 ;
      RECT 470.065 -35.545 480.215 2.225 ;
      RECT 451.385 -34.825 465.315 2.225 ;
      RECT 455.165 -35.545 465.315 2.225 ;
      RECT 436.485 -34.825 450.415 2.225 ;
      RECT 440.265 -35.545 450.415 2.225 ;
      RECT 421.585 -34.825 435.515 2.225 ;
      RECT 425.365 -35.545 435.515 2.225 ;
      RECT 406.685 -34.825 420.615 2.225 ;
      RECT 410.465 -35.545 420.615 2.225 ;
      RECT 391.785 -34.825 405.715 2.225 ;
      RECT 395.565 -35.545 405.715 2.225 ;
      RECT 376.885 -34.825 390.815 2.225 ;
      RECT 380.665 -35.545 390.815 2.225 ;
      RECT 361.985 -34.825 375.915 2.225 ;
      RECT 365.765 -35.545 375.915 2.225 ;
      RECT 347.085 -34.825 361.015 2.225 ;
      RECT 350.865 -35.545 361.015 2.225 ;
      RECT 332.185 -34.825 346.115 2.225 ;
      RECT 335.965 -35.545 346.115 2.225 ;
      RECT 317.285 -34.825 331.215 2.225 ;
      RECT 321.065 -35.545 331.215 2.225 ;
      RECT 302.385 -34.825 316.315 2.225 ;
      RECT 306.165 -35.545 316.315 2.225 ;
      RECT 287.485 -34.825 301.415 2.225 ;
      RECT 291.265 -35.545 301.415 2.225 ;
      RECT 272.585 -34.825 286.515 2.225 ;
      RECT 276.365 -35.545 286.515 2.225 ;
      RECT 257.685 -34.825 271.615 2.225 ;
      RECT 261.465 -35.545 271.615 2.225 ;
      RECT 242.785 -34.825 256.715 2.225 ;
      RECT 246.565 -35.545 256.715 2.225 ;
      RECT 227.885 -34.825 241.815 2.225 ;
      RECT 231.665 -35.545 241.815 2.225 ;
      RECT 212.985 -34.825 226.915 2.225 ;
      RECT 216.765 -35.545 226.915 2.225 ;
      RECT 198.085 -34.825 212.015 2.225 ;
      RECT 201.865 -35.545 212.015 2.225 ;
      RECT 183.185 -34.825 197.115 2.225 ;
      RECT 186.965 -35.545 197.115 2.225 ;
      RECT 168.285 -34.825 182.215 2.225 ;
      RECT 172.065 -35.545 182.215 2.225 ;
      RECT 153.385 -34.825 167.315 2.225 ;
      RECT 157.165 -35.545 167.315 2.225 ;
      RECT 138.485 -34.825 152.415 2.225 ;
      RECT 142.265 -35.545 152.415 2.225 ;
      RECT 123.585 -34.825 137.515 2.225 ;
      RECT 127.365 -35.545 137.515 2.225 ;
      RECT 108.685 -34.825 122.615 2.225 ;
      RECT 112.465 -35.545 122.615 2.225 ;
      RECT 93.785 -34.825 107.715 2.225 ;
      RECT 97.565 -35.545 107.715 2.225 ;
      RECT 78.885 -34.825 92.815 2.225 ;
      RECT 82.665 -35.545 92.815 2.225 ;
      RECT 63.985 -34.825 77.915 2.225 ;
      RECT 67.765 -35.545 77.915 2.225 ;
      RECT 49.085 -34.825 63.015 2.225 ;
      RECT 52.865 -35.545 63.015 2.225 ;
      RECT 34.185 -34.825 48.115 2.225 ;
      RECT 37.965 -35.545 48.115 2.225 ;
      RECT 19.285 -34.825 33.215 2.225 ;
      RECT 23.065 -35.545 33.215 2.225 ;
      RECT 6.905 -34.825 18.315 2.225 ;
      RECT 8.165 -35.545 18.315 2.225 ;
      RECT -1.525 -35.545 5.935 2.225 ;
      RECT 945.605 -35.545 945.895 2.225 ;
      RECT 930.705 -35.545 930.995 2.225 ;
      RECT 929.445 -35.545 929.735 2.225 ;
      RECT 928.185 -35.545 928.475 2.225 ;
      RECT 915.805 -35.545 916.095 2.225 ;
      RECT 914.545 -35.545 914.835 2.225 ;
      RECT 913.285 -35.545 913.575 2.225 ;
      RECT 900.905 -35.545 901.195 2.225 ;
      RECT 899.645 -35.545 899.935 2.225 ;
      RECT 898.385 -35.545 898.675 2.225 ;
      RECT 886.005 -35.545 886.295 2.225 ;
      RECT 884.745 -35.545 885.035 2.225 ;
      RECT 883.485 -35.545 883.775 2.225 ;
      RECT 871.105 -35.545 871.395 2.225 ;
      RECT 869.845 -35.545 870.135 2.225 ;
      RECT 868.585 -35.545 868.875 2.225 ;
      RECT 856.205 -35.545 856.495 2.225 ;
      RECT 854.945 -35.545 855.235 2.225 ;
      RECT 853.685 -35.545 853.975 2.225 ;
      RECT 841.305 -35.545 841.595 2.225 ;
      RECT 840.045 -35.545 840.335 2.225 ;
      RECT 838.785 -35.545 839.075 2.225 ;
      RECT 826.405 -35.545 826.695 2.225 ;
      RECT 825.145 -35.545 825.435 2.225 ;
      RECT 823.885 -35.545 824.175 2.225 ;
      RECT 811.505 -35.545 811.795 2.225 ;
      RECT 810.245 -35.545 810.535 2.225 ;
      RECT 808.985 -35.545 809.275 2.225 ;
      RECT 796.605 -35.545 796.895 2.225 ;
      RECT 795.345 -35.545 795.635 2.225 ;
      RECT 794.085 -35.545 794.375 2.225 ;
      RECT 781.705 -35.545 781.995 2.225 ;
      RECT 780.445 -35.545 780.735 2.225 ;
      RECT 779.185 -35.545 779.475 2.225 ;
      RECT 766.805 -35.545 767.095 2.225 ;
      RECT 765.545 -35.545 765.835 2.225 ;
      RECT 764.285 -35.545 764.575 2.225 ;
      RECT 751.905 -35.545 752.195 2.225 ;
      RECT 750.645 -35.545 750.935 2.225 ;
      RECT 749.385 -35.545 749.675 2.225 ;
      RECT 737.005 -35.545 737.295 2.225 ;
      RECT 735.745 -35.545 736.035 2.225 ;
      RECT 734.485 -35.545 734.775 2.225 ;
      RECT 722.105 -35.545 722.395 2.225 ;
      RECT 720.845 -35.545 721.135 2.225 ;
      RECT 719.585 -35.545 719.875 2.225 ;
      RECT 707.205 -35.545 707.495 2.225 ;
      RECT 705.945 -35.545 706.235 2.225 ;
      RECT 704.685 -35.545 704.975 2.225 ;
      RECT 692.305 -35.545 692.595 2.225 ;
      RECT 691.045 -35.545 691.335 2.225 ;
      RECT 689.785 -35.545 690.075 2.225 ;
      RECT 677.405 -35.545 677.695 2.225 ;
      RECT 676.145 -35.545 676.435 2.225 ;
      RECT 674.885 -35.545 675.175 2.225 ;
      RECT 662.505 -35.545 662.795 2.225 ;
      RECT 661.245 -35.545 661.535 2.225 ;
      RECT 659.985 -35.545 660.275 2.225 ;
      RECT 647.605 -35.545 647.895 2.225 ;
      RECT 646.345 -35.545 646.635 2.225 ;
      RECT 645.085 -35.545 645.375 2.225 ;
      RECT 632.705 -35.545 632.995 2.225 ;
      RECT 631.445 -35.545 631.735 2.225 ;
      RECT 630.185 -35.545 630.475 2.225 ;
      RECT 617.805 -35.545 618.095 2.225 ;
      RECT 616.545 -35.545 616.835 2.225 ;
      RECT 615.285 -35.545 615.575 2.225 ;
      RECT 602.905 -35.545 603.195 2.225 ;
      RECT 601.645 -35.545 601.935 2.225 ;
      RECT 600.385 -35.545 600.675 2.225 ;
      RECT 588.005 -35.545 588.295 2.225 ;
      RECT 586.745 -35.545 587.035 2.225 ;
      RECT 585.485 -35.545 585.775 2.225 ;
      RECT 573.105 -35.545 573.395 2.225 ;
      RECT 571.845 -35.545 572.135 2.225 ;
      RECT 570.585 -35.545 570.875 2.225 ;
      RECT 558.205 -35.545 558.495 2.225 ;
      RECT 556.945 -35.545 557.235 2.225 ;
      RECT 555.685 -35.545 555.975 2.225 ;
      RECT 543.305 -35.545 543.595 2.225 ;
      RECT 542.045 -35.545 542.335 2.225 ;
      RECT 540.785 -35.545 541.075 2.225 ;
      RECT 528.405 -35.545 528.695 2.225 ;
      RECT 527.145 -35.545 527.435 2.225 ;
      RECT 525.885 -35.545 526.175 2.225 ;
      RECT 513.505 -35.545 513.795 2.225 ;
      RECT 512.245 -35.545 512.535 2.225 ;
      RECT 510.985 -35.545 511.275 2.225 ;
      RECT 498.605 -35.545 498.895 2.225 ;
      RECT 497.345 -35.545 497.635 2.225 ;
      RECT 496.085 -35.545 496.375 2.225 ;
      RECT 483.705 -35.545 483.995 2.225 ;
      RECT 482.445 -35.545 482.735 2.225 ;
      RECT 481.185 -35.545 481.475 2.225 ;
      RECT 468.805 -35.545 469.095 2.225 ;
      RECT 467.545 -35.545 467.835 2.225 ;
      RECT 466.285 -35.545 466.575 2.225 ;
      RECT 453.905 -35.545 454.195 2.225 ;
      RECT 452.645 -35.545 452.935 2.225 ;
      RECT 451.385 -35.545 451.675 2.225 ;
      RECT 439.005 -35.545 439.295 2.225 ;
      RECT 437.745 -35.545 438.035 2.225 ;
      RECT 436.485 -35.545 436.775 2.225 ;
      RECT 424.105 -35.545 424.395 2.225 ;
      RECT 422.845 -35.545 423.135 2.225 ;
      RECT 421.585 -35.545 421.875 2.225 ;
      RECT 409.205 -35.545 409.495 2.225 ;
      RECT 407.945 -35.545 408.235 2.225 ;
      RECT 406.685 -35.545 406.975 2.225 ;
      RECT 394.305 -35.545 394.595 2.225 ;
      RECT 393.045 -35.545 393.335 2.225 ;
      RECT 391.785 -35.545 392.075 2.225 ;
      RECT 379.405 -35.545 379.695 2.225 ;
      RECT 378.145 -35.545 378.435 2.225 ;
      RECT 376.885 -35.545 377.175 2.225 ;
      RECT 364.505 -35.545 364.795 2.225 ;
      RECT 363.245 -35.545 363.535 2.225 ;
      RECT 361.985 -35.545 362.275 2.225 ;
      RECT 349.605 -35.545 349.895 2.225 ;
      RECT 348.345 -35.545 348.635 2.225 ;
      RECT 347.085 -35.545 347.375 2.225 ;
      RECT 334.705 -35.545 334.995 2.225 ;
      RECT 333.445 -35.545 333.735 2.225 ;
      RECT 332.185 -35.545 332.475 2.225 ;
      RECT 319.805 -35.545 320.095 2.225 ;
      RECT 318.545 -35.545 318.835 2.225 ;
      RECT 317.285 -35.545 317.575 2.225 ;
      RECT 304.905 -35.545 305.195 2.225 ;
      RECT 303.645 -35.545 303.935 2.225 ;
      RECT 302.385 -35.545 302.675 2.225 ;
      RECT 290.005 -35.545 290.295 2.225 ;
      RECT 288.745 -35.545 289.035 2.225 ;
      RECT 287.485 -35.545 287.775 2.225 ;
      RECT 275.105 -35.545 275.395 2.225 ;
      RECT 273.845 -35.545 274.135 2.225 ;
      RECT 272.585 -35.545 272.875 2.225 ;
      RECT 260.205 -35.545 260.495 2.225 ;
      RECT 258.945 -35.545 259.235 2.225 ;
      RECT 257.685 -35.545 257.975 2.225 ;
      RECT 245.305 -35.545 245.595 2.225 ;
      RECT 244.045 -35.545 244.335 2.225 ;
      RECT 242.785 -35.545 243.075 2.225 ;
      RECT 230.405 -35.545 230.695 2.225 ;
      RECT 229.145 -35.545 229.435 2.225 ;
      RECT 227.885 -35.545 228.175 2.225 ;
      RECT 215.505 -35.545 215.795 2.225 ;
      RECT 214.245 -35.545 214.535 2.225 ;
      RECT 212.985 -35.545 213.275 2.225 ;
      RECT 200.605 -35.545 200.895 2.225 ;
      RECT 199.345 -35.545 199.635 2.225 ;
      RECT 198.085 -35.545 198.375 2.225 ;
      RECT 185.705 -35.545 185.995 2.225 ;
      RECT 184.445 -35.545 184.735 2.225 ;
      RECT 183.185 -35.545 183.475 2.225 ;
      RECT 170.805 -35.545 171.095 2.225 ;
      RECT 169.545 -35.545 169.835 2.225 ;
      RECT 168.285 -35.545 168.575 2.225 ;
      RECT 155.905 -35.545 156.195 2.225 ;
      RECT 154.645 -35.545 154.935 2.225 ;
      RECT 153.385 -35.545 153.675 2.225 ;
      RECT 141.005 -35.545 141.295 2.225 ;
      RECT 139.745 -35.545 140.035 2.225 ;
      RECT 138.485 -35.545 138.775 2.225 ;
      RECT 126.105 -35.545 126.395 2.225 ;
      RECT 124.845 -35.545 125.135 2.225 ;
      RECT 123.585 -35.545 123.875 2.225 ;
      RECT 111.205 -35.545 111.495 2.225 ;
      RECT 109.945 -35.545 110.235 2.225 ;
      RECT 108.685 -35.545 108.975 2.225 ;
      RECT 96.305 -35.545 96.595 2.225 ;
      RECT 95.045 -35.545 95.335 2.225 ;
      RECT 93.785 -35.545 94.075 2.225 ;
      RECT 81.405 -35.545 81.695 2.225 ;
      RECT 80.145 -35.545 80.435 2.225 ;
      RECT 78.885 -35.545 79.175 2.225 ;
      RECT 66.505 -35.545 66.795 2.225 ;
      RECT 65.245 -35.545 65.535 2.225 ;
      RECT 63.985 -35.545 64.275 2.225 ;
      RECT 51.605 -35.545 51.895 2.225 ;
      RECT 50.345 -35.545 50.635 2.225 ;
      RECT 49.085 -35.545 49.375 2.225 ;
      RECT 36.705 -35.545 36.995 2.225 ;
      RECT 35.445 -35.545 35.735 2.225 ;
      RECT 34.185 -35.545 34.475 2.225 ;
      RECT 21.805 -35.545 22.095 2.225 ;
      RECT 20.545 -35.545 20.835 2.225 ;
      RECT 19.285 -35.545 19.575 2.225 ;
      RECT 6.905 -35.545 7.195 2.225 ;
    LAYER met3 SPACING 0.3 ;
      RECT -0.54 -24.725 954.04 -24.395 ;
      RECT -0.54 -22.025 954.04 -21.695 ;
      RECT 944.955 -35.475 948.435 -35.145 ;
      RECT 942.435 -22.875 944.025 -22.545 ;
      RECT 941.805 -23.505 942.765 -23.175 ;
      RECT 927.535 -35.475 934.165 -35.145 ;
      RECT 928.795 -29.805 934.165 -29.475 ;
      RECT 931.315 -26.655 934.165 -26.325 ;
      RECT 927.535 -27.915 930.385 -27.585 ;
      RECT 927.535 -23.505 929.755 -23.175 ;
      RECT 927.535 -22.875 929.125 -22.545 ;
      RECT 926.905 -29.805 927.865 -29.475 ;
      RECT 912.635 -35.475 919.265 -35.145 ;
      RECT 913.895 -29.805 919.265 -29.475 ;
      RECT 916.415 -26.655 919.265 -26.325 ;
      RECT 912.635 -27.915 915.485 -27.585 ;
      RECT 912.635 -23.505 914.855 -23.175 ;
      RECT 912.635 -22.875 914.225 -22.545 ;
      RECT 912.005 -29.805 912.965 -29.475 ;
      RECT 897.735 -35.475 904.365 -35.145 ;
      RECT 898.995 -29.805 904.365 -29.475 ;
      RECT 901.515 -26.655 904.365 -26.325 ;
      RECT 897.735 -27.915 900.585 -27.585 ;
      RECT 897.735 -23.505 899.955 -23.175 ;
      RECT 897.735 -22.875 899.325 -22.545 ;
      RECT 897.105 -29.805 898.065 -29.475 ;
      RECT 882.835 -35.475 889.465 -35.145 ;
      RECT 884.095 -29.805 889.465 -29.475 ;
      RECT 886.615 -26.655 889.465 -26.325 ;
      RECT 882.835 -27.915 885.685 -27.585 ;
      RECT 882.835 -23.505 885.055 -23.175 ;
      RECT 882.835 -22.875 884.425 -22.545 ;
      RECT 882.205 -29.805 883.165 -29.475 ;
      RECT 867.935 -35.475 874.565 -35.145 ;
      RECT 869.195 -29.805 874.565 -29.475 ;
      RECT 871.715 -26.655 874.565 -26.325 ;
      RECT 867.935 -27.915 870.785 -27.585 ;
      RECT 867.935 -23.505 870.155 -23.175 ;
      RECT 867.935 -22.875 869.525 -22.545 ;
      RECT 867.305 -29.805 868.265 -29.475 ;
      RECT 853.035 -35.475 859.665 -35.145 ;
      RECT 854.295 -29.805 859.665 -29.475 ;
      RECT 856.815 -26.655 859.665 -26.325 ;
      RECT 853.035 -27.915 855.885 -27.585 ;
      RECT 853.035 -23.505 855.255 -23.175 ;
      RECT 853.035 -22.875 854.625 -22.545 ;
      RECT 852.405 -29.805 853.365 -29.475 ;
      RECT 838.135 -35.475 844.765 -35.145 ;
      RECT 839.395 -29.805 844.765 -29.475 ;
      RECT 841.915 -26.655 844.765 -26.325 ;
      RECT 838.135 -27.915 840.985 -27.585 ;
      RECT 838.135 -23.505 840.355 -23.175 ;
      RECT 838.135 -22.875 839.725 -22.545 ;
      RECT 837.505 -29.805 838.465 -29.475 ;
      RECT 823.235 -35.475 829.865 -35.145 ;
      RECT 824.495 -29.805 829.865 -29.475 ;
      RECT 827.015 -26.655 829.865 -26.325 ;
      RECT 823.235 -27.915 826.085 -27.585 ;
      RECT 823.235 -23.505 825.455 -23.175 ;
      RECT 823.235 -22.875 824.825 -22.545 ;
      RECT 822.605 -29.805 823.565 -29.475 ;
      RECT 808.335 -35.475 814.965 -35.145 ;
      RECT 809.595 -29.805 814.965 -29.475 ;
      RECT 812.115 -26.655 814.965 -26.325 ;
      RECT 808.335 -27.915 811.185 -27.585 ;
      RECT 808.335 -23.505 810.555 -23.175 ;
      RECT 808.335 -22.875 809.925 -22.545 ;
      RECT 807.705 -29.805 808.665 -29.475 ;
      RECT 793.435 -35.475 800.065 -35.145 ;
      RECT 794.695 -29.805 800.065 -29.475 ;
      RECT 797.215 -26.655 800.065 -26.325 ;
      RECT 793.435 -27.915 796.285 -27.585 ;
      RECT 793.435 -23.505 795.655 -23.175 ;
      RECT 793.435 -22.875 795.025 -22.545 ;
      RECT 792.805 -29.805 793.765 -29.475 ;
      RECT 778.535 -35.475 785.165 -35.145 ;
      RECT 779.795 -29.805 785.165 -29.475 ;
      RECT 782.315 -26.655 785.165 -26.325 ;
      RECT 778.535 -27.915 781.385 -27.585 ;
      RECT 778.535 -23.505 780.755 -23.175 ;
      RECT 778.535 -22.875 780.125 -22.545 ;
      RECT 777.905 -29.805 778.865 -29.475 ;
      RECT 763.635 -35.475 770.265 -35.145 ;
      RECT 764.895 -29.805 770.265 -29.475 ;
      RECT 767.415 -26.655 770.265 -26.325 ;
      RECT 763.635 -27.915 766.485 -27.585 ;
      RECT 763.635 -23.505 765.855 -23.175 ;
      RECT 763.635 -22.875 765.225 -22.545 ;
      RECT 763.005 -29.805 763.965 -29.475 ;
      RECT 748.735 -35.475 755.365 -35.145 ;
      RECT 749.995 -29.805 755.365 -29.475 ;
      RECT 752.515 -26.655 755.365 -26.325 ;
      RECT 748.735 -27.915 751.585 -27.585 ;
      RECT 748.735 -23.505 750.955 -23.175 ;
      RECT 748.735 -22.875 750.325 -22.545 ;
      RECT 748.105 -29.805 749.065 -29.475 ;
      RECT 733.835 -35.475 740.465 -35.145 ;
      RECT 735.095 -29.805 740.465 -29.475 ;
      RECT 737.615 -26.655 740.465 -26.325 ;
      RECT 733.835 -27.915 736.685 -27.585 ;
      RECT 733.835 -23.505 736.055 -23.175 ;
      RECT 733.835 -22.875 735.425 -22.545 ;
      RECT 733.205 -29.805 734.165 -29.475 ;
      RECT 718.935 -35.475 725.565 -35.145 ;
      RECT 720.195 -29.805 725.565 -29.475 ;
      RECT 722.715 -26.655 725.565 -26.325 ;
      RECT 718.935 -27.915 721.785 -27.585 ;
      RECT 718.935 -23.505 721.155 -23.175 ;
      RECT 718.935 -22.875 720.525 -22.545 ;
      RECT 718.305 -29.805 719.265 -29.475 ;
      RECT 704.035 -35.475 710.665 -35.145 ;
      RECT 705.295 -29.805 710.665 -29.475 ;
      RECT 707.815 -26.655 710.665 -26.325 ;
      RECT 704.035 -27.915 706.885 -27.585 ;
      RECT 704.035 -23.505 706.255 -23.175 ;
      RECT 704.035 -22.875 705.625 -22.545 ;
      RECT 703.405 -29.805 704.365 -29.475 ;
      RECT 689.135 -35.475 695.765 -35.145 ;
      RECT 690.395 -29.805 695.765 -29.475 ;
      RECT 692.915 -26.655 695.765 -26.325 ;
      RECT 689.135 -27.915 691.985 -27.585 ;
      RECT 689.135 -23.505 691.355 -23.175 ;
      RECT 689.135 -22.875 690.725 -22.545 ;
      RECT 688.505 -29.805 689.465 -29.475 ;
      RECT 674.235 -35.475 680.865 -35.145 ;
      RECT 675.495 -29.805 680.865 -29.475 ;
      RECT 678.015 -26.655 680.865 -26.325 ;
      RECT 674.235 -27.915 677.085 -27.585 ;
      RECT 674.235 -23.505 676.455 -23.175 ;
      RECT 674.235 -22.875 675.825 -22.545 ;
      RECT 673.605 -29.805 674.565 -29.475 ;
      RECT 659.335 -35.475 665.965 -35.145 ;
      RECT 660.595 -29.805 665.965 -29.475 ;
      RECT 663.115 -26.655 665.965 -26.325 ;
      RECT 659.335 -27.915 662.185 -27.585 ;
      RECT 659.335 -23.505 661.555 -23.175 ;
      RECT 659.335 -22.875 660.925 -22.545 ;
      RECT 658.705 -29.805 659.665 -29.475 ;
      RECT 644.435 -35.475 651.065 -35.145 ;
      RECT 645.695 -29.805 651.065 -29.475 ;
      RECT 648.215 -26.655 651.065 -26.325 ;
      RECT 644.435 -27.915 647.285 -27.585 ;
      RECT 644.435 -23.505 646.655 -23.175 ;
      RECT 644.435 -22.875 646.025 -22.545 ;
      RECT 643.805 -29.805 644.765 -29.475 ;
      RECT 629.535 -35.475 636.165 -35.145 ;
      RECT 630.795 -29.805 636.165 -29.475 ;
      RECT 633.315 -26.655 636.165 -26.325 ;
      RECT 629.535 -27.915 632.385 -27.585 ;
      RECT 629.535 -23.505 631.755 -23.175 ;
      RECT 629.535 -22.875 631.125 -22.545 ;
      RECT 628.905 -29.805 629.865 -29.475 ;
      RECT 614.635 -35.475 621.265 -35.145 ;
      RECT 615.895 -29.805 621.265 -29.475 ;
      RECT 618.415 -26.655 621.265 -26.325 ;
      RECT 614.635 -27.915 617.485 -27.585 ;
      RECT 614.635 -23.505 616.855 -23.175 ;
      RECT 614.635 -22.875 616.225 -22.545 ;
      RECT 614.005 -29.805 614.965 -29.475 ;
      RECT 599.735 -35.475 606.365 -35.145 ;
      RECT 600.995 -29.805 606.365 -29.475 ;
      RECT 603.515 -26.655 606.365 -26.325 ;
      RECT 599.735 -27.915 602.585 -27.585 ;
      RECT 599.735 -23.505 601.955 -23.175 ;
      RECT 599.735 -22.875 601.325 -22.545 ;
      RECT 599.105 -29.805 600.065 -29.475 ;
      RECT 584.835 -35.475 591.465 -35.145 ;
      RECT 586.095 -29.805 591.465 -29.475 ;
      RECT 588.615 -26.655 591.465 -26.325 ;
      RECT 584.835 -27.915 587.685 -27.585 ;
      RECT 584.835 -23.505 587.055 -23.175 ;
      RECT 584.835 -22.875 586.425 -22.545 ;
      RECT 584.205 -29.805 585.165 -29.475 ;
      RECT 569.935 -35.475 576.565 -35.145 ;
      RECT 571.195 -29.805 576.565 -29.475 ;
      RECT 573.715 -26.655 576.565 -26.325 ;
      RECT 569.935 -27.915 572.785 -27.585 ;
      RECT 569.935 -23.505 572.155 -23.175 ;
      RECT 569.935 -22.875 571.525 -22.545 ;
      RECT 569.305 -29.805 570.265 -29.475 ;
      RECT 555.035 -35.475 561.665 -35.145 ;
      RECT 556.295 -29.805 561.665 -29.475 ;
      RECT 558.815 -26.655 561.665 -26.325 ;
      RECT 555.035 -27.915 557.885 -27.585 ;
      RECT 555.035 -23.505 557.255 -23.175 ;
      RECT 555.035 -22.875 556.625 -22.545 ;
      RECT 554.405 -29.805 555.365 -29.475 ;
      RECT 540.135 -35.475 546.765 -35.145 ;
      RECT 541.395 -29.805 546.765 -29.475 ;
      RECT 543.915 -26.655 546.765 -26.325 ;
      RECT 540.135 -27.915 542.985 -27.585 ;
      RECT 540.135 -23.505 542.355 -23.175 ;
      RECT 540.135 -22.875 541.725 -22.545 ;
      RECT 539.505 -29.805 540.465 -29.475 ;
      RECT 525.235 -35.475 531.865 -35.145 ;
      RECT 526.495 -29.805 531.865 -29.475 ;
      RECT 529.015 -26.655 531.865 -26.325 ;
      RECT 525.235 -27.915 528.085 -27.585 ;
      RECT 525.235 -23.505 527.455 -23.175 ;
      RECT 525.235 -22.875 526.825 -22.545 ;
      RECT 524.605 -29.805 525.565 -29.475 ;
      RECT 510.335 -35.475 516.965 -35.145 ;
      RECT 511.595 -29.805 516.965 -29.475 ;
      RECT 514.115 -26.655 516.965 -26.325 ;
      RECT 510.335 -27.915 513.185 -27.585 ;
      RECT 510.335 -23.505 512.555 -23.175 ;
      RECT 510.335 -22.875 511.925 -22.545 ;
      RECT 509.705 -29.805 510.665 -29.475 ;
      RECT 495.435 -35.475 502.065 -35.145 ;
      RECT 496.695 -29.805 502.065 -29.475 ;
      RECT 499.215 -26.655 502.065 -26.325 ;
      RECT 495.435 -27.915 498.285 -27.585 ;
      RECT 495.435 -23.505 497.655 -23.175 ;
      RECT 495.435 -22.875 497.025 -22.545 ;
      RECT 494.805 -29.805 495.765 -29.475 ;
      RECT 480.535 -35.475 487.165 -35.145 ;
      RECT 481.795 -29.805 487.165 -29.475 ;
      RECT 484.315 -26.655 487.165 -26.325 ;
      RECT 480.535 -27.915 483.385 -27.585 ;
      RECT 480.535 -23.505 482.755 -23.175 ;
      RECT 480.535 -22.875 482.125 -22.545 ;
      RECT 479.905 -29.805 480.865 -29.475 ;
      RECT 465.635 -35.475 472.265 -35.145 ;
      RECT 466.895 -29.805 472.265 -29.475 ;
      RECT 469.415 -26.655 472.265 -26.325 ;
      RECT 465.635 -27.915 468.485 -27.585 ;
      RECT 465.635 -23.505 467.855 -23.175 ;
      RECT 465.635 -22.875 467.225 -22.545 ;
      RECT 465.005 -29.805 465.965 -29.475 ;
      RECT 450.735 -35.475 457.365 -35.145 ;
      RECT 451.995 -29.805 457.365 -29.475 ;
      RECT 454.515 -26.655 457.365 -26.325 ;
      RECT 450.735 -27.915 453.585 -27.585 ;
      RECT 450.735 -23.505 452.955 -23.175 ;
      RECT 450.735 -22.875 452.325 -22.545 ;
      RECT 450.105 -29.805 451.065 -29.475 ;
      RECT 435.835 -35.475 442.465 -35.145 ;
      RECT 437.095 -29.805 442.465 -29.475 ;
      RECT 439.615 -26.655 442.465 -26.325 ;
      RECT 435.835 -27.915 438.685 -27.585 ;
      RECT 435.835 -23.505 438.055 -23.175 ;
      RECT 435.835 -22.875 437.425 -22.545 ;
      RECT 435.205 -29.805 436.165 -29.475 ;
      RECT 420.935 -35.475 427.565 -35.145 ;
      RECT 422.195 -29.805 427.565 -29.475 ;
      RECT 424.715 -26.655 427.565 -26.325 ;
      RECT 420.935 -27.915 423.785 -27.585 ;
      RECT 420.935 -23.505 423.155 -23.175 ;
      RECT 420.935 -22.875 422.525 -22.545 ;
      RECT 420.305 -29.805 421.265 -29.475 ;
      RECT 406.035 -35.475 412.665 -35.145 ;
      RECT 407.295 -29.805 412.665 -29.475 ;
      RECT 409.815 -26.655 412.665 -26.325 ;
      RECT 406.035 -27.915 408.885 -27.585 ;
      RECT 406.035 -23.505 408.255 -23.175 ;
      RECT 406.035 -22.875 407.625 -22.545 ;
      RECT 405.405 -29.805 406.365 -29.475 ;
      RECT 391.135 -35.475 397.765 -35.145 ;
      RECT 392.395 -29.805 397.765 -29.475 ;
      RECT 394.915 -26.655 397.765 -26.325 ;
      RECT 391.135 -27.915 393.985 -27.585 ;
      RECT 391.135 -23.505 393.355 -23.175 ;
      RECT 391.135 -22.875 392.725 -22.545 ;
      RECT 390.505 -29.805 391.465 -29.475 ;
      RECT 376.235 -35.475 382.865 -35.145 ;
      RECT 377.495 -29.805 382.865 -29.475 ;
      RECT 380.015 -26.655 382.865 -26.325 ;
      RECT 376.235 -27.915 379.085 -27.585 ;
      RECT 376.235 -23.505 378.455 -23.175 ;
      RECT 376.235 -22.875 377.825 -22.545 ;
      RECT 375.605 -29.805 376.565 -29.475 ;
      RECT 361.335 -35.475 367.965 -35.145 ;
      RECT 362.595 -29.805 367.965 -29.475 ;
      RECT 365.115 -26.655 367.965 -26.325 ;
      RECT 361.335 -27.915 364.185 -27.585 ;
      RECT 361.335 -23.505 363.555 -23.175 ;
      RECT 361.335 -22.875 362.925 -22.545 ;
      RECT 360.705 -29.805 361.665 -29.475 ;
      RECT 346.435 -35.475 353.065 -35.145 ;
      RECT 347.695 -29.805 353.065 -29.475 ;
      RECT 350.215 -26.655 353.065 -26.325 ;
      RECT 346.435 -27.915 349.285 -27.585 ;
      RECT 346.435 -23.505 348.655 -23.175 ;
      RECT 346.435 -22.875 348.025 -22.545 ;
      RECT 345.805 -29.805 346.765 -29.475 ;
      RECT 331.535 -35.475 338.165 -35.145 ;
      RECT 332.795 -29.805 338.165 -29.475 ;
      RECT 335.315 -26.655 338.165 -26.325 ;
      RECT 331.535 -27.915 334.385 -27.585 ;
      RECT 331.535 -23.505 333.755 -23.175 ;
      RECT 331.535 -22.875 333.125 -22.545 ;
      RECT 330.905 -29.805 331.865 -29.475 ;
      RECT 316.635 -35.475 323.265 -35.145 ;
      RECT 317.895 -29.805 323.265 -29.475 ;
      RECT 320.415 -26.655 323.265 -26.325 ;
      RECT 316.635 -27.915 319.485 -27.585 ;
      RECT 316.635 -23.505 318.855 -23.175 ;
      RECT 316.635 -22.875 318.225 -22.545 ;
      RECT 316.005 -29.805 316.965 -29.475 ;
      RECT 301.735 -35.475 308.365 -35.145 ;
      RECT 302.995 -29.805 308.365 -29.475 ;
      RECT 305.515 -26.655 308.365 -26.325 ;
      RECT 301.735 -27.915 304.585 -27.585 ;
      RECT 301.735 -23.505 303.955 -23.175 ;
      RECT 301.735 -22.875 303.325 -22.545 ;
      RECT 301.105 -29.805 302.065 -29.475 ;
      RECT 286.835 -35.475 293.465 -35.145 ;
      RECT 288.095 -29.805 293.465 -29.475 ;
      RECT 290.615 -26.655 293.465 -26.325 ;
      RECT 286.835 -27.915 289.685 -27.585 ;
      RECT 286.835 -23.505 289.055 -23.175 ;
      RECT 286.835 -22.875 288.425 -22.545 ;
      RECT 286.205 -29.805 287.165 -29.475 ;
      RECT 271.935 -35.475 278.565 -35.145 ;
      RECT 273.195 -29.805 278.565 -29.475 ;
      RECT 275.715 -26.655 278.565 -26.325 ;
      RECT 271.935 -27.915 274.785 -27.585 ;
      RECT 271.935 -23.505 274.155 -23.175 ;
      RECT 271.935 -22.875 273.525 -22.545 ;
      RECT 271.305 -29.805 272.265 -29.475 ;
      RECT 257.035 -35.475 263.665 -35.145 ;
      RECT 258.295 -29.805 263.665 -29.475 ;
      RECT 260.815 -26.655 263.665 -26.325 ;
      RECT 257.035 -27.915 259.885 -27.585 ;
      RECT 257.035 -23.505 259.255 -23.175 ;
      RECT 257.035 -22.875 258.625 -22.545 ;
      RECT 256.405 -29.805 257.365 -29.475 ;
      RECT 242.135 -35.475 248.765 -35.145 ;
      RECT 243.395 -29.805 248.765 -29.475 ;
      RECT 245.915 -26.655 248.765 -26.325 ;
      RECT 242.135 -27.915 244.985 -27.585 ;
      RECT 242.135 -23.505 244.355 -23.175 ;
      RECT 242.135 -22.875 243.725 -22.545 ;
      RECT 241.505 -29.805 242.465 -29.475 ;
      RECT 227.235 -35.475 233.865 -35.145 ;
      RECT 228.495 -29.805 233.865 -29.475 ;
      RECT 231.015 -26.655 233.865 -26.325 ;
      RECT 227.235 -27.915 230.085 -27.585 ;
      RECT 227.235 -23.505 229.455 -23.175 ;
      RECT 227.235 -22.875 228.825 -22.545 ;
      RECT 226.605 -29.805 227.565 -29.475 ;
      RECT 212.335 -35.475 218.965 -35.145 ;
      RECT 213.595 -29.805 218.965 -29.475 ;
      RECT 216.115 -26.655 218.965 -26.325 ;
      RECT 212.335 -27.915 215.185 -27.585 ;
      RECT 212.335 -23.505 214.555 -23.175 ;
      RECT 212.335 -22.875 213.925 -22.545 ;
      RECT 211.705 -29.805 212.665 -29.475 ;
      RECT 197.435 -35.475 204.065 -35.145 ;
      RECT 198.695 -29.805 204.065 -29.475 ;
      RECT 201.215 -26.655 204.065 -26.325 ;
      RECT 197.435 -27.915 200.285 -27.585 ;
      RECT 197.435 -23.505 199.655 -23.175 ;
      RECT 197.435 -22.875 199.025 -22.545 ;
      RECT 196.805 -29.805 197.765 -29.475 ;
      RECT 182.535 -35.475 189.165 -35.145 ;
      RECT 183.795 -29.805 189.165 -29.475 ;
      RECT 186.315 -26.655 189.165 -26.325 ;
      RECT 182.535 -27.915 185.385 -27.585 ;
      RECT 182.535 -23.505 184.755 -23.175 ;
      RECT 182.535 -22.875 184.125 -22.545 ;
      RECT 181.905 -29.805 182.865 -29.475 ;
      RECT 167.635 -35.475 174.265 -35.145 ;
      RECT 168.895 -29.805 174.265 -29.475 ;
      RECT 171.415 -26.655 174.265 -26.325 ;
      RECT 167.635 -27.915 170.485 -27.585 ;
      RECT 167.635 -23.505 169.855 -23.175 ;
      RECT 167.635 -22.875 169.225 -22.545 ;
      RECT 167.005 -29.805 167.965 -29.475 ;
      RECT 152.735 -35.475 159.365 -35.145 ;
      RECT 153.995 -29.805 159.365 -29.475 ;
      RECT 156.515 -26.655 159.365 -26.325 ;
      RECT 152.735 -27.915 155.585 -27.585 ;
      RECT 152.735 -23.505 154.955 -23.175 ;
      RECT 152.735 -22.875 154.325 -22.545 ;
      RECT 152.105 -29.805 153.065 -29.475 ;
      RECT 137.835 -35.475 144.465 -35.145 ;
      RECT 139.095 -29.805 144.465 -29.475 ;
      RECT 141.615 -26.655 144.465 -26.325 ;
      RECT 137.835 -27.915 140.685 -27.585 ;
      RECT 137.835 -23.505 140.055 -23.175 ;
      RECT 137.835 -22.875 139.425 -22.545 ;
      RECT 137.205 -29.805 138.165 -29.475 ;
      RECT 122.935 -35.475 129.565 -35.145 ;
      RECT 124.195 -29.805 129.565 -29.475 ;
      RECT 126.715 -26.655 129.565 -26.325 ;
      RECT 122.935 -27.915 125.785 -27.585 ;
      RECT 122.935 -23.505 125.155 -23.175 ;
      RECT 122.935 -22.875 124.525 -22.545 ;
      RECT 122.305 -29.805 123.265 -29.475 ;
      RECT 108.035 -35.475 114.665 -35.145 ;
      RECT 109.295 -29.805 114.665 -29.475 ;
      RECT 111.815 -26.655 114.665 -26.325 ;
      RECT 108.035 -27.915 110.885 -27.585 ;
      RECT 108.035 -23.505 110.255 -23.175 ;
      RECT 108.035 -22.875 109.625 -22.545 ;
      RECT 107.405 -29.805 108.365 -29.475 ;
      RECT 93.135 -35.475 99.765 -35.145 ;
      RECT 94.395 -29.805 99.765 -29.475 ;
      RECT 96.915 -26.655 99.765 -26.325 ;
      RECT 93.135 -27.915 95.985 -27.585 ;
      RECT 93.135 -23.505 95.355 -23.175 ;
      RECT 93.135 -22.875 94.725 -22.545 ;
      RECT 92.505 -29.805 93.465 -29.475 ;
      RECT 78.235 -35.475 84.865 -35.145 ;
      RECT 79.495 -29.805 84.865 -29.475 ;
      RECT 82.015 -26.655 84.865 -26.325 ;
      RECT 78.235 -27.915 81.085 -27.585 ;
      RECT 78.235 -23.505 80.455 -23.175 ;
      RECT 78.235 -22.875 79.825 -22.545 ;
      RECT 77.605 -29.805 78.565 -29.475 ;
      RECT 63.335 -35.475 69.965 -35.145 ;
      RECT 64.595 -29.805 69.965 -29.475 ;
      RECT 67.115 -26.655 69.965 -26.325 ;
      RECT 63.335 -27.915 66.185 -27.585 ;
      RECT 63.335 -23.505 65.555 -23.175 ;
      RECT 63.335 -22.875 64.925 -22.545 ;
      RECT 62.705 -29.805 63.665 -29.475 ;
      RECT 48.435 -35.475 55.065 -35.145 ;
      RECT 49.695 -29.805 55.065 -29.475 ;
      RECT 52.215 -26.655 55.065 -26.325 ;
      RECT 48.435 -27.915 51.285 -27.585 ;
      RECT 48.435 -23.505 50.655 -23.175 ;
      RECT 48.435 -22.875 50.025 -22.545 ;
      RECT 47.805 -29.805 48.765 -29.475 ;
      RECT 33.535 -35.475 40.165 -35.145 ;
      RECT 34.795 -29.805 40.165 -29.475 ;
      RECT 37.315 -26.655 40.165 -26.325 ;
      RECT 33.535 -27.915 36.385 -27.585 ;
      RECT 33.535 -23.505 35.755 -23.175 ;
      RECT 33.535 -22.875 35.125 -22.545 ;
      RECT 32.905 -29.805 33.865 -29.475 ;
      RECT 18.635 -35.475 25.265 -35.145 ;
      RECT 19.895 -29.805 25.265 -29.475 ;
      RECT 22.415 -26.655 25.265 -26.325 ;
      RECT 18.635 -27.915 21.485 -27.585 ;
      RECT 18.635 -23.505 20.855 -23.175 ;
      RECT 18.635 -22.875 20.225 -22.545 ;
      RECT 18.005 -29.805 18.965 -29.475 ;
      RECT 6.255 -35.475 9.735 -35.145 ;
      RECT 3.735 -23.505 5.955 -23.175 ;
      RECT 3.735 -22.875 5.325 -22.545 ;
  END
END tdc_64

END LIBRARY
